-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to 24575) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80d6",
     9 => x"f4080b0b",
    10 => x"80d6f808",
    11 => x"0b0b80d6",
    12 => x"fc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"d6fc0c0b",
    16 => x"0b80d6f8",
    17 => x"0c0b0b80",
    18 => x"d6f40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80cfa8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80d6f470",
    57 => x"81c9b027",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c5188f7",
    62 => x"04820b0b",
    63 => x"0b80d2e0",
    64 => x"0c800b80",
    65 => x"d78c0c80",
    66 => x"0b80d784",
    67 => x"0c800b80",
    68 => x"d7880c04",
    69 => x"02fc050d",
    70 => x"f880518f",
    71 => x"0b80d784",
    72 => x"0c9f0b80",
    73 => x"d7880ca0",
    74 => x"71708105",
    75 => x"533480d7",
    76 => x"8808ff05",
    77 => x"80d7880c",
    78 => x"80d78808",
    79 => x"8025e838",
    80 => x"80d78408",
    81 => x"ff0580d7",
    82 => x"840c80d7",
    83 => x"84088025",
    84 => x"d038800b",
    85 => x"80d7880c",
    86 => x"800b80d7",
    87 => x"840c0284",
    88 => x"050d0402",
    89 => x"f0050df8",
    90 => x"8053f8a0",
    91 => x"5483bf52",
    92 => x"73708105",
    93 => x"55335170",
    94 => x"73708105",
    95 => x"5534ff12",
    96 => x"52718025",
    97 => x"eb38fbc0",
    98 => x"539f52a0",
    99 => x"73708105",
   100 => x"5534ff12",
   101 => x"52718025",
   102 => x"f2380290",
   103 => x"050d0402",
   104 => x"f4050d74",
   105 => x"538e0b80",
   106 => x"d7840825",
   107 => x"913882e3",
   108 => x"2d80d784",
   109 => x"08ff0580",
   110 => x"d7840c83",
   111 => x"a50480d7",
   112 => x"840880d7",
   113 => x"88085351",
   114 => x"728a2e09",
   115 => x"8106be38",
   116 => x"7151719f",
   117 => x"24a43880",
   118 => x"d78408a0",
   119 => x"2911f880",
   120 => x"115151a0",
   121 => x"713480d7",
   122 => x"88088105",
   123 => x"80d7880c",
   124 => x"80d78808",
   125 => x"519f7125",
   126 => x"de38800b",
   127 => x"80d7880c",
   128 => x"80d78408",
   129 => x"810580d7",
   130 => x"840c84a3",
   131 => x"0470a029",
   132 => x"12f88011",
   133 => x"51517271",
   134 => x"3480d788",
   135 => x"08810580",
   136 => x"d7880c80",
   137 => x"d78808a0",
   138 => x"2e098106",
   139 => x"9138800b",
   140 => x"80d7880c",
   141 => x"80d78408",
   142 => x"810580d7",
   143 => x"840c028c",
   144 => x"050d0402",
   145 => x"e8050d77",
   146 => x"79565688",
   147 => x"0bfc1677",
   148 => x"712c8f06",
   149 => x"54525480",
   150 => x"53727225",
   151 => x"95387153",
   152 => x"fbe01451",
   153 => x"87713481",
   154 => x"14ff1454",
   155 => x"5472f138",
   156 => x"7153f915",
   157 => x"76712c87",
   158 => x"06535171",
   159 => x"802e8b38",
   160 => x"fbe01451",
   161 => x"71713481",
   162 => x"1454728e",
   163 => x"2495388f",
   164 => x"733153fb",
   165 => x"e01451a0",
   166 => x"71348114",
   167 => x"ff145454",
   168 => x"72f13802",
   169 => x"98050d04",
   170 => x"02f4050d",
   171 => x"800b80d7",
   172 => x"8c0cf68c",
   173 => x"08f69008",
   174 => x"71882c72",
   175 => x"81ff0653",
   176 => x"54545171",
   177 => x"71258738",
   178 => x"820b80d7",
   179 => x"8c0c7288",
   180 => x"2c7381ff",
   181 => x"06525271",
   182 => x"71258b38",
   183 => x"80d78c08",
   184 => x"840780d7",
   185 => x"8c0c820b",
   186 => x"0b0b80d2",
   187 => x"e00c830b",
   188 => x"f6880cfc",
   189 => x"0880d78c",
   190 => x"08515174",
   191 => x"802e8538",
   192 => x"70810751",
   193 => x"70f6940c",
   194 => x"feb80bf6",
   195 => x"800cff9c",
   196 => x"0bf6840c",
   197 => x"028c050d",
   198 => x"0402f405",
   199 => x"0d745372",
   200 => x"70810554",
   201 => x"80f52d52",
   202 => x"71802e89",
   203 => x"38715183",
   204 => x"9f2d869f",
   205 => x"04810b80",
   206 => x"d6f40c02",
   207 => x"8c050d04",
   208 => x"02f0050d",
   209 => x"76537552",
   210 => x"80d4a80b",
   211 => x"80f52d51",
   212 => x"80cba72d",
   213 => x"80d6f408",
   214 => x"5480d6f4",
   215 => x"08802e88",
   216 => x"3880d388",
   217 => x"5186ec04",
   218 => x"80d48451",
   219 => x"90cd2d73",
   220 => x"80d6f40c",
   221 => x"0290050d",
   222 => x"0402fc05",
   223 => x"0d800b80",
   224 => x"d4a80b81",
   225 => x"b72d86c0",
   226 => x"5180c498",
   227 => x"2d725180",
   228 => x"c3f32d02",
   229 => x"84050d04",
   230 => x"02fc050d",
   231 => x"810b80d4",
   232 => x"a80b81b7",
   233 => x"2d86c051",
   234 => x"80c4982d",
   235 => x"725180c3",
   236 => x"f32d0284",
   237 => x"050d0402",
   238 => x"f4050d74",
   239 => x"53805180",
   240 => x"d48008a7",
   241 => x"24a03870",
   242 => x"52711351",
   243 => x"807181b7",
   244 => x"2d811252",
   245 => x"83ff7225",
   246 => x"f03880d4",
   247 => x"80088105",
   248 => x"80d4800c",
   249 => x"81517080",
   250 => x"d6f40c02",
   251 => x"8c050d04",
   252 => x"02c8050d",
   253 => x"800b80d0",
   254 => x"ec53029c",
   255 => x"05705356",
   256 => x"5680cdd5",
   257 => x"2d745202",
   258 => x"a8055488",
   259 => x"9b047552",
   260 => x"81167552",
   261 => x"5680cea8",
   262 => x"2d745273",
   263 => x"5180cdd5",
   264 => x"2d80d0f4",
   265 => x"52735180",
   266 => x"cdf72d73",
   267 => x"51b9d22d",
   268 => x"80d6f408",
   269 => x"d93880d0",
   270 => x"fc518699",
   271 => x"2d735186",
   272 => x"992d80d1",
   273 => x"ec518699",
   274 => x"2d800b80",
   275 => x"d4800cb2",
   276 => x"80805387",
   277 => x"b7527351",
   278 => x"80c4c12d",
   279 => x"80d6f408",
   280 => x"802e8838",
   281 => x"80d38851",
   282 => x"88ef0480",
   283 => x"d4845190",
   284 => x"cd2d02b8",
   285 => x"050d0402",
   286 => x"f4050df0",
   287 => x"08810652",
   288 => x"8ae42d8c",
   289 => x"da2d8f92",
   290 => x"2d9de62d",
   291 => x"81f92d71",
   292 => x"8538850b",
   293 => x"ec0c8ef7",
   294 => x"2d8a892d",
   295 => x"82942d81",
   296 => x"5185a82d",
   297 => x"840bec0c",
   298 => x"80d18c51",
   299 => x"86992da1",
   300 => x"8c2d80d6",
   301 => x"f408802e",
   302 => x"b73880cc",
   303 => x"8d2d80d2",
   304 => x"e45190cd",
   305 => x"2d805185",
   306 => x"a82d840b",
   307 => x"ec0c8b9b",
   308 => x"2d90e02d",
   309 => x"80d6f408",
   310 => x"5280cadc",
   311 => x"2d80d4fc",
   312 => x"08fc0c86",
   313 => x"53718338",
   314 => x"845372ec",
   315 => x"0c89ce04",
   316 => x"800b80d6",
   317 => x"f40c028c",
   318 => x"050d0480",
   319 => x"0bffb00c",
   320 => x"04ffb008",
   321 => x"80d6f40c",
   322 => x"04810bff",
   323 => x"b00c0402",
   324 => x"f8050d89",
   325 => x"fb2d8a81",
   326 => x"2d80d6f4",
   327 => x"0880d790",
   328 => x"0880d6f4",
   329 => x"083280d7",
   330 => x"900c80d6",
   331 => x"f4088106",
   332 => x"52527080",
   333 => x"2e8d3880",
   334 => x"d4ac0851",
   335 => x"70802e83",
   336 => x"38702d71",
   337 => x"812a7081",
   338 => x"06515170",
   339 => x"802e8d38",
   340 => x"80d4b008",
   341 => x"5170802e",
   342 => x"8338702d",
   343 => x"8a892d02",
   344 => x"88050d04",
   345 => x"02fc050d",
   346 => x"80d4ac51",
   347 => x"80717084",
   348 => x"05530c80",
   349 => x"710c0284",
   350 => x"050d0402",
   351 => x"fc050d72",
   352 => x"8a8f0b98",
   353 => x"0c517081",
   354 => x"248c3870",
   355 => x"842980d4",
   356 => x"ac057471",
   357 => x"0c510284",
   358 => x"050d0402",
   359 => x"f4050d80",
   360 => x"d794518e",
   361 => x"812d80d6",
   362 => x"f4085280",
   363 => x"d6f40880",
   364 => x"2e819d38",
   365 => x"8cbe0480",
   366 => x"d6f40881",
   367 => x"f02e0981",
   368 => x"068a3881",
   369 => x"0b80d4f4",
   370 => x"0c8cbe04",
   371 => x"80d6f408",
   372 => x"81e02e09",
   373 => x"81068a38",
   374 => x"810b80d4",
   375 => x"f80c8cbe",
   376 => x"0480d6f4",
   377 => x"085280d4",
   378 => x"f808802e",
   379 => x"893880d6",
   380 => x"f4088180",
   381 => x"05527184",
   382 => x"2c728f06",
   383 => x"535380d4",
   384 => x"f408802e",
   385 => x"9a387284",
   386 => x"2980d4b4",
   387 => x"05721381",
   388 => x"712b7009",
   389 => x"73080673",
   390 => x"0c515353",
   391 => x"8cb20472",
   392 => x"842980d4",
   393 => x"b4057213",
   394 => x"83712b72",
   395 => x"0807720c",
   396 => x"5353800b",
   397 => x"80d4f80c",
   398 => x"800b80d4",
   399 => x"f40c80d7",
   400 => x"94518dbc",
   401 => x"2d80d6f4",
   402 => x"08ff24fe",
   403 => x"ea388052",
   404 => x"7180d6f4",
   405 => x"0c028c05",
   406 => x"0d0402f8",
   407 => x"050d80d4",
   408 => x"b4528f51",
   409 => x"80727084",
   410 => x"05540cff",
   411 => x"11517080",
   412 => x"25f23802",
   413 => x"88050d04",
   414 => x"02f0050d",
   415 => x"7570822c",
   416 => x"fc0680d4",
   417 => x"b4117210",
   418 => x"9e067108",
   419 => x"70722a82",
   420 => x"732b7009",
   421 => x"7306750c",
   422 => x"53830680",
   423 => x"d6f40c57",
   424 => x"53515351",
   425 => x"0290050d",
   426 => x"0402fc05",
   427 => x"0d725180",
   428 => x"710c800b",
   429 => x"84120c02",
   430 => x"84050d04",
   431 => x"02f0050d",
   432 => x"75700884",
   433 => x"12085353",
   434 => x"53ff5471",
   435 => x"712ea838",
   436 => x"89fb2d84",
   437 => x"13087084",
   438 => x"29148811",
   439 => x"70087081",
   440 => x"ff068418",
   441 => x"08811187",
   442 => x"06841a0c",
   443 => x"53515551",
   444 => x"51518a89",
   445 => x"2d715473",
   446 => x"80d6f40c",
   447 => x"0290050d",
   448 => x"0402f405",
   449 => x"0d747008",
   450 => x"84120853",
   451 => x"53537072",
   452 => x"248f3872",
   453 => x"08841408",
   454 => x"71713152",
   455 => x"52528eae",
   456 => x"04720884",
   457 => x"14087171",
   458 => x"31880552",
   459 => x"52527180",
   460 => x"d6f40c02",
   461 => x"8c050d04",
   462 => x"02f8050d",
   463 => x"e008708b",
   464 => x"2a708106",
   465 => x"51525270",
   466 => x"802ea138",
   467 => x"80d79408",
   468 => x"70842980",
   469 => x"d79c0573",
   470 => x"81ff0671",
   471 => x"0c515180",
   472 => x"d7940881",
   473 => x"11870680",
   474 => x"d7940c51",
   475 => x"800b80d7",
   476 => x"bc0c0288",
   477 => x"050d0402",
   478 => x"f8050d80",
   479 => x"d794518d",
   480 => x"a92d8cda",
   481 => x"2d8eb852",
   482 => x"80518afb",
   483 => x"2d028805",
   484 => x"0d04800b",
   485 => x"80d5800c",
   486 => x"81c60b80",
   487 => x"d4fc0c04",
   488 => x"80d7c008",
   489 => x"80d6f40c",
   490 => x"0402fc05",
   491 => x"0d8fb304",
   492 => x"8b9b2d87",
   493 => x"518cf82d",
   494 => x"80d6f408",
   495 => x"f33880da",
   496 => x"518cf82d",
   497 => x"80d6f408",
   498 => x"e73880d6",
   499 => x"f40880d5",
   500 => x"800c80d6",
   501 => x"f4085185",
   502 => x"a82d0284",
   503 => x"050d0402",
   504 => x"f4050d80",
   505 => x"d7c00853",
   506 => x"82942d80",
   507 => x"0b80d7c4",
   508 => x"0c720880",
   509 => x"2e80d138",
   510 => x"820b80d7",
   511 => x"880c80d7",
   512 => x"c4088f06",
   513 => x"80d7840c",
   514 => x"7208812e",
   515 => x"098106a1",
   516 => x"3880d4fc",
   517 => x"08881408",
   518 => x"2c708106",
   519 => x"51527180",
   520 => x"2e883880",
   521 => x"d1a45190",
   522 => x"ae0480d1",
   523 => x"a8518699",
   524 => x"2d841308",
   525 => x"5186992d",
   526 => x"80d7c408",
   527 => x"810580d7",
   528 => x"c40c8c13",
   529 => x"538ff104",
   530 => x"028c050d",
   531 => x"047180d7",
   532 => x"c00c8fdf",
   533 => x"2d80d7c4",
   534 => x"08ff0580",
   535 => x"d7c80c04",
   536 => x"02e8050d",
   537 => x"80d7c008",
   538 => x"80d7cc08",
   539 => x"56568751",
   540 => x"8cf82d80",
   541 => x"d6f40881",
   542 => x"2a708106",
   543 => x"51527180",
   544 => x"2eac3891",
   545 => x"89048b9b",
   546 => x"2d87518c",
   547 => x"f82d80d6",
   548 => x"f408f338",
   549 => x"80d58008",
   550 => x"81327080",
   551 => x"d5800c51",
   552 => x"85a82d80",
   553 => x"d5800880",
   554 => x"2e84388c",
   555 => x"da2d80d5",
   556 => x"80087054",
   557 => x"5271802e",
   558 => x"84a63881",
   559 => x"f5518cf8",
   560 => x"2d80d6f4",
   561 => x"08812a70",
   562 => x"81065152",
   563 => x"71802eb3",
   564 => x"3880d7c8",
   565 => x"08527180",
   566 => x"2e8a38ff",
   567 => x"1280d7c8",
   568 => x"0c928304",
   569 => x"80d7c408",
   570 => x"1080d7c4",
   571 => x"08057084",
   572 => x"29175152",
   573 => x"88120880",
   574 => x"2e8938ff",
   575 => x"51881208",
   576 => x"52712d81",
   577 => x"f2518cf8",
   578 => x"2d80d6f4",
   579 => x"08812a70",
   580 => x"81065152",
   581 => x"71802eb4",
   582 => x"3880d7c4",
   583 => x"08ff1180",
   584 => x"d7c80856",
   585 => x"53537372",
   586 => x"258a3881",
   587 => x"1480d7c8",
   588 => x"0c92cc04",
   589 => x"72101370",
   590 => x"84291751",
   591 => x"52881208",
   592 => x"802e8938",
   593 => x"fe518812",
   594 => x"0852712d",
   595 => x"81fd518c",
   596 => x"f82d80d6",
   597 => x"f408812a",
   598 => x"70810651",
   599 => x"5271802e",
   600 => x"b13880d7",
   601 => x"c808802e",
   602 => x"8a38800b",
   603 => x"80d7c80c",
   604 => x"93920480",
   605 => x"d7c40810",
   606 => x"80d7c408",
   607 => x"05708429",
   608 => x"17515288",
   609 => x"1208802e",
   610 => x"8938fd51",
   611 => x"88120852",
   612 => x"712d81fa",
   613 => x"518cf82d",
   614 => x"80d6f408",
   615 => x"812a7081",
   616 => x"06515271",
   617 => x"802eb138",
   618 => x"80d7c408",
   619 => x"ff115452",
   620 => x"80d7c808",
   621 => x"73258938",
   622 => x"7280d7c8",
   623 => x"0c93d804",
   624 => x"71101270",
   625 => x"84291751",
   626 => x"52881208",
   627 => x"802e8938",
   628 => x"fc518812",
   629 => x"0852712d",
   630 => x"80d7c808",
   631 => x"70535473",
   632 => x"802e8738",
   633 => x"ff145493",
   634 => x"df04820b",
   635 => x"80d7880c",
   636 => x"718f0680",
   637 => x"d7840c80",
   638 => x"da518cf8",
   639 => x"2d80d6f4",
   640 => x"08812a70",
   641 => x"81065152",
   642 => x"71802e81",
   643 => x"8a3880d7",
   644 => x"c00880d7",
   645 => x"c8085553",
   646 => x"73802e8a",
   647 => x"388c13ff",
   648 => x"15555394",
   649 => x"98047208",
   650 => x"5271822e",
   651 => x"a1387182",
   652 => x"26893871",
   653 => x"812ea538",
   654 => x"95970471",
   655 => x"842e0981",
   656 => x"0680d438",
   657 => x"88130851",
   658 => x"90cd2d95",
   659 => x"970480d7",
   660 => x"c8085188",
   661 => x"13085271",
   662 => x"2d959704",
   663 => x"810b8814",
   664 => x"082b80d4",
   665 => x"fc083280",
   666 => x"d4fc0c8f",
   667 => x"df2d9597",
   668 => x"04740880",
   669 => x"2ea43874",
   670 => x"08518cf8",
   671 => x"2d80d6f4",
   672 => x"08810652",
   673 => x"71802e8c",
   674 => x"3880d7c8",
   675 => x"08518415",
   676 => x"0852712d",
   677 => x"88155574",
   678 => x"d8388054",
   679 => x"800b80d7",
   680 => x"880c738f",
   681 => x"0680d784",
   682 => x"0ca05273",
   683 => x"80d7c808",
   684 => x"2e098106",
   685 => x"993880d7",
   686 => x"c408ff05",
   687 => x"74327009",
   688 => x"81057072",
   689 => x"079f2a91",
   690 => x"71315151",
   691 => x"53537151",
   692 => x"839f2d81",
   693 => x"14548e74",
   694 => x"25c23880",
   695 => x"d5800853",
   696 => x"7280d6f4",
   697 => x"0c029805",
   698 => x"0d0402f4",
   699 => x"050dd452",
   700 => x"81ff720c",
   701 => x"71085381",
   702 => x"ff720c72",
   703 => x"882b83fe",
   704 => x"80067208",
   705 => x"7081ff06",
   706 => x"51525381",
   707 => x"ff720c72",
   708 => x"7107882b",
   709 => x"72087081",
   710 => x"ff065152",
   711 => x"5381ff72",
   712 => x"0c727107",
   713 => x"882b7208",
   714 => x"7081ff06",
   715 => x"720780d6",
   716 => x"f40c5253",
   717 => x"028c050d",
   718 => x"0402f405",
   719 => x"0d747671",
   720 => x"81ff06d4",
   721 => x"0c535380",
   722 => x"d7d00885",
   723 => x"3871892b",
   724 => x"5271982a",
   725 => x"d40c7190",
   726 => x"2a7081ff",
   727 => x"06d40c51",
   728 => x"71882a70",
   729 => x"81ff06d4",
   730 => x"0c517181",
   731 => x"ff06d40c",
   732 => x"72902a70",
   733 => x"81ff06d4",
   734 => x"0c51d408",
   735 => x"7081ff06",
   736 => x"515182b8",
   737 => x"bf527081",
   738 => x"ff2e0981",
   739 => x"06943881",
   740 => x"ff0bd40c",
   741 => x"d4087081",
   742 => x"ff06ff14",
   743 => x"54515171",
   744 => x"e5387080",
   745 => x"d6f40c02",
   746 => x"8c050d04",
   747 => x"02fc050d",
   748 => x"81c75181",
   749 => x"ff0bd40c",
   750 => x"ff115170",
   751 => x"8025f438",
   752 => x"0284050d",
   753 => x"0402f405",
   754 => x"0d81ff0b",
   755 => x"d40c9353",
   756 => x"805287fc",
   757 => x"80c15196",
   758 => x"b92d80d6",
   759 => x"f4088b38",
   760 => x"81ff0bd4",
   761 => x"0c815397",
   762 => x"f30497ac",
   763 => x"2dff1353",
   764 => x"72de3872",
   765 => x"80d6f40c",
   766 => x"028c050d",
   767 => x"0402ec05",
   768 => x"0d810b80",
   769 => x"d7d00c84",
   770 => x"54d00870",
   771 => x"8f2a7081",
   772 => x"06515153",
   773 => x"72f33872",
   774 => x"d00c97ac",
   775 => x"2d80d1ac",
   776 => x"5186992d",
   777 => x"d008708f",
   778 => x"2a708106",
   779 => x"51515372",
   780 => x"f338810b",
   781 => x"d00cb153",
   782 => x"805284d4",
   783 => x"80c05196",
   784 => x"b92d80d6",
   785 => x"f408812e",
   786 => x"93387282",
   787 => x"2ebf38ff",
   788 => x"135372e4",
   789 => x"38ff1454",
   790 => x"73ffae38",
   791 => x"97ac2d83",
   792 => x"aa52849c",
   793 => x"80c85196",
   794 => x"b92d80d6",
   795 => x"f408812e",
   796 => x"09810693",
   797 => x"3895ea2d",
   798 => x"80d6f408",
   799 => x"83ffff06",
   800 => x"537283aa",
   801 => x"2e9f3897",
   802 => x"c52d99a0",
   803 => x"0480d1b8",
   804 => x"5186992d",
   805 => x"80539af5",
   806 => x"0480d1d0",
   807 => x"5186992d",
   808 => x"80549ac6",
   809 => x"0481ff0b",
   810 => x"d40cb154",
   811 => x"97ac2d8f",
   812 => x"cf538052",
   813 => x"87fc80f7",
   814 => x"5196b92d",
   815 => x"80d6f408",
   816 => x"5580d6f4",
   817 => x"08812e09",
   818 => x"81069c38",
   819 => x"81ff0bd4",
   820 => x"0c820a52",
   821 => x"849c80e9",
   822 => x"5196b92d",
   823 => x"80d6f408",
   824 => x"802e8d38",
   825 => x"97ac2dff",
   826 => x"135372c6",
   827 => x"389ab904",
   828 => x"81ff0bd4",
   829 => x"0c80d6f4",
   830 => x"085287fc",
   831 => x"80fa5196",
   832 => x"b92d80d6",
   833 => x"f408b238",
   834 => x"81ff0bd4",
   835 => x"0cd40853",
   836 => x"81ff0bd4",
   837 => x"0c81ff0b",
   838 => x"d40c81ff",
   839 => x"0bd40c81",
   840 => x"ff0bd40c",
   841 => x"72862a70",
   842 => x"81067656",
   843 => x"51537296",
   844 => x"3880d6f4",
   845 => x"08549ac6",
   846 => x"0473822e",
   847 => x"fedb38ff",
   848 => x"145473fe",
   849 => x"e7387380",
   850 => x"d7d00c73",
   851 => x"8b388152",
   852 => x"87fc80d0",
   853 => x"5196b92d",
   854 => x"81ff0bd4",
   855 => x"0cd00870",
   856 => x"8f2a7081",
   857 => x"06515153",
   858 => x"72f33872",
   859 => x"d00c81ff",
   860 => x"0bd40c81",
   861 => x"537280d6",
   862 => x"f40c0294",
   863 => x"050d0402",
   864 => x"e8050d78",
   865 => x"5681ff0b",
   866 => x"d40cd008",
   867 => x"708f2a70",
   868 => x"81065151",
   869 => x"5372f338",
   870 => x"82810bd0",
   871 => x"0c81ff0b",
   872 => x"d40c7752",
   873 => x"87fc80d8",
   874 => x"5196b92d",
   875 => x"80d6f408",
   876 => x"802e8d38",
   877 => x"80d1e051",
   878 => x"86992d81",
   879 => x"539cb804",
   880 => x"81ff0bd4",
   881 => x"0c81fe0b",
   882 => x"d40c80ff",
   883 => x"55757084",
   884 => x"05570870",
   885 => x"982ad40c",
   886 => x"70902c70",
   887 => x"81ff06d4",
   888 => x"0c547088",
   889 => x"2c7081ff",
   890 => x"06d40c54",
   891 => x"7081ff06",
   892 => x"d40c54ff",
   893 => x"15557480",
   894 => x"25d33881",
   895 => x"ff0bd40c",
   896 => x"81ff0bd4",
   897 => x"0c81ff0b",
   898 => x"d40c868d",
   899 => x"a05481ff",
   900 => x"0bd40cd4",
   901 => x"0881ff06",
   902 => x"55748738",
   903 => x"ff145473",
   904 => x"ed3881ff",
   905 => x"0bd40cd0",
   906 => x"08708f2a",
   907 => x"70810651",
   908 => x"515372f3",
   909 => x"3872d00c",
   910 => x"7280d6f4",
   911 => x"0c029805",
   912 => x"0d0402e8",
   913 => x"050d7855",
   914 => x"805681ff",
   915 => x"0bd40cd0",
   916 => x"08708f2a",
   917 => x"70810651",
   918 => x"515372f3",
   919 => x"3882810b",
   920 => x"d00c81ff",
   921 => x"0bd40c77",
   922 => x"5287fc80",
   923 => x"d15196b9",
   924 => x"2d80dbc6",
   925 => x"df5480d6",
   926 => x"f408802e",
   927 => x"8b3880d1",
   928 => x"f0518699",
   929 => x"2d9ddc04",
   930 => x"81ff0bd4",
   931 => x"0cd40870",
   932 => x"81ff0651",
   933 => x"537281fe",
   934 => x"2e098106",
   935 => x"9e3880ff",
   936 => x"5395ea2d",
   937 => x"80d6f408",
   938 => x"75708405",
   939 => x"570cff13",
   940 => x"53728025",
   941 => x"ec388156",
   942 => x"9dc104ff",
   943 => x"145473c8",
   944 => x"3881ff0b",
   945 => x"d40c81ff",
   946 => x"0bd40cd0",
   947 => x"08708f2a",
   948 => x"70810651",
   949 => x"515372f3",
   950 => x"3872d00c",
   951 => x"7580d6f4",
   952 => x"0c029805",
   953 => x"0d04800b",
   954 => x"80dde80c",
   955 => x"800b80dd",
   956 => x"ec0c800b",
   957 => x"80dde00c",
   958 => x"800b80dd",
   959 => x"f00c800b",
   960 => x"80ddf40c",
   961 => x"800b80dd",
   962 => x"f80c800b",
   963 => x"80ddfc0c",
   964 => x"800b80de",
   965 => x"800c800b",
   966 => x"80de840c",
   967 => x"800b80dd",
   968 => x"d80c800b",
   969 => x"80dddc0c",
   970 => x"800b80de",
   971 => x"880c800b",
   972 => x"80de8c0c",
   973 => x"800b80de",
   974 => x"900b818a",
   975 => x"2d820b80",
   976 => x"d58c0c80",
   977 => x"0b80de94",
   978 => x"0c800b80",
   979 => x"de980c80",
   980 => x"0b80de9c",
   981 => x"0c800b80",
   982 => x"dea00c80",
   983 => x"0b80dde4",
   984 => x"0c800b80",
   985 => x"d5840c04",
   986 => x"02e8050d",
   987 => x"77797b58",
   988 => x"55558053",
   989 => x"727625a3",
   990 => x"38747081",
   991 => x"055680f5",
   992 => x"2d747081",
   993 => x"055680f5",
   994 => x"2d525271",
   995 => x"712e8638",
   996 => x"81519f9d",
   997 => x"04811353",
   998 => x"9ef40480",
   999 => x"517080d6",
  1000 => x"f40c0298",
  1001 => x"050d0402",
  1002 => x"f8050d73",
  1003 => x"5280dde0",
  1004 => x"08802e94",
  1005 => x"3871822b",
  1006 => x"83fc0680",
  1007 => x"dea41108",
  1008 => x"5252be8a",
  1009 => x"2d9fd904",
  1010 => x"711083fe",
  1011 => x"0680dea4",
  1012 => x"1180e02d",
  1013 => x"5252beb5",
  1014 => x"2d028805",
  1015 => x"0d0402ec",
  1016 => x"050d7655",
  1017 => x"74802e80",
  1018 => x"c5389a15",
  1019 => x"80e02d51",
  1020 => x"beb52d80",
  1021 => x"d6f40880",
  1022 => x"d6f40880",
  1023 => x"de980c80",
  1024 => x"d6f40854",
  1025 => x"5480dde0",
  1026 => x"08802e9a",
  1027 => x"38941580",
  1028 => x"e02d51be",
  1029 => x"b52d80d6",
  1030 => x"f408902b",
  1031 => x"83fff00a",
  1032 => x"06707507",
  1033 => x"51537280",
  1034 => x"de980ca0",
  1035 => x"b3047480",
  1036 => x"de980c80",
  1037 => x"de980853",
  1038 => x"72802e9d",
  1039 => x"3880ddd8",
  1040 => x"08fe1471",
  1041 => x"2980ddf4",
  1042 => x"080580de",
  1043 => x"9c0c7084",
  1044 => x"2b80dde4",
  1045 => x"0c54a187",
  1046 => x"0480ddf8",
  1047 => x"0880de98",
  1048 => x"0c80ddfc",
  1049 => x"0880de9c",
  1050 => x"0c80dde0",
  1051 => x"08802e8b",
  1052 => x"3880ddd8",
  1053 => x"08842b53",
  1054 => x"a1820480",
  1055 => x"de800884",
  1056 => x"2b537280",
  1057 => x"dde40c02",
  1058 => x"94050d04",
  1059 => x"02d8050d",
  1060 => x"800b80dd",
  1061 => x"e00c8454",
  1062 => x"97fd2d80",
  1063 => x"d6f40880",
  1064 => x"2e973880",
  1065 => x"d7d45280",
  1066 => x"519cc22d",
  1067 => x"80d6f408",
  1068 => x"802e8638",
  1069 => x"fe54a1c1",
  1070 => x"04ff1454",
  1071 => x"738024d8",
  1072 => x"38738d38",
  1073 => x"80d28051",
  1074 => x"86992d73",
  1075 => x"55a8da04",
  1076 => x"800b80de",
  1077 => x"940c810b",
  1078 => x"80dea00c",
  1079 => x"885380d2",
  1080 => x"945280d8",
  1081 => x"8a519ee8",
  1082 => x"2d80d6f4",
  1083 => x"08893880",
  1084 => x"d6f40880",
  1085 => x"dea00c88",
  1086 => x"5380d2a0",
  1087 => x"5280d8a6",
  1088 => x"519ee82d",
  1089 => x"80d6f408",
  1090 => x"893880d6",
  1091 => x"f40880de",
  1092 => x"a00c80de",
  1093 => x"a008802e",
  1094 => x"818c3880",
  1095 => x"db9a0b80",
  1096 => x"f52d80db",
  1097 => x"9b0b80f5",
  1098 => x"2d71982b",
  1099 => x"71902b07",
  1100 => x"80db9c0b",
  1101 => x"80f52d70",
  1102 => x"882b7207",
  1103 => x"80db9d0b",
  1104 => x"80f52d71",
  1105 => x"077080de",
  1106 => x"940c80db",
  1107 => x"d20b80f5",
  1108 => x"2d80dbd3",
  1109 => x"0b80f52d",
  1110 => x"71882b07",
  1111 => x"575f5152",
  1112 => x"5a565755",
  1113 => x"7481abaa",
  1114 => x"2e098106",
  1115 => x"91387351",
  1116 => x"be8a2d80",
  1117 => x"d6f40880",
  1118 => x"de940ca3",
  1119 => x"8c047482",
  1120 => x"d4d52e88",
  1121 => x"3880d2ac",
  1122 => x"51a3db04",
  1123 => x"80d7d452",
  1124 => x"80de9408",
  1125 => x"519cc22d",
  1126 => x"80d6f408",
  1127 => x"5580d6f4",
  1128 => x"08802e85",
  1129 => x"b5388853",
  1130 => x"80d2a052",
  1131 => x"80d8a651",
  1132 => x"9ee82d80",
  1133 => x"d6f4088a",
  1134 => x"38810b80",
  1135 => x"dde00ca3",
  1136 => x"e1048853",
  1137 => x"80d29452",
  1138 => x"80d88a51",
  1139 => x"9ee82d80",
  1140 => x"d6f40880",
  1141 => x"2e8b3880",
  1142 => x"d2c05186",
  1143 => x"992da4c0",
  1144 => x"0480dbd2",
  1145 => x"0b80f52d",
  1146 => x"547380d5",
  1147 => x"2e098106",
  1148 => x"80ce3880",
  1149 => x"dbd30b80",
  1150 => x"f52d5473",
  1151 => x"81aa2e09",
  1152 => x"8106bd38",
  1153 => x"800b80d7",
  1154 => x"d40b80f5",
  1155 => x"2d565474",
  1156 => x"81e92e83",
  1157 => x"38815474",
  1158 => x"81eb2e8c",
  1159 => x"38805573",
  1160 => x"752e0981",
  1161 => x"0684b338",
  1162 => x"80d7df0b",
  1163 => x"80f52d56",
  1164 => x"758e3880",
  1165 => x"d7e00b80",
  1166 => x"f52d5473",
  1167 => x"822e8638",
  1168 => x"8055a8da",
  1169 => x"0480d7e1",
  1170 => x"0b80f52d",
  1171 => x"7080ddd8",
  1172 => x"0cff0570",
  1173 => x"80dddc0c",
  1174 => x"55817680",
  1175 => x"de880c70",
  1176 => x"76065557",
  1177 => x"73802e97",
  1178 => x"38747656",
  1179 => x"58811577",
  1180 => x"10707a06",
  1181 => x"56585573",
  1182 => x"f4387480",
  1183 => x"de880c80",
  1184 => x"d7e20b80",
  1185 => x"f52d80d7",
  1186 => x"e30b80f5",
  1187 => x"2d5680de",
  1188 => x"94080575",
  1189 => x"82802905",
  1190 => x"7080ddf0",
  1191 => x"0c80d7e4",
  1192 => x"0b80f52d",
  1193 => x"7080de84",
  1194 => x"0c80dde0",
  1195 => x"08595758",
  1196 => x"76802e82",
  1197 => x"c6388853",
  1198 => x"80d2a052",
  1199 => x"80d8a651",
  1200 => x"9ee82d80",
  1201 => x"5580d6f4",
  1202 => x"08752e09",
  1203 => x"8106838a",
  1204 => x"3880ddd8",
  1205 => x"0870842b",
  1206 => x"80dde40c",
  1207 => x"7080de80",
  1208 => x"0c80d7f9",
  1209 => x"0b80f52d",
  1210 => x"80d7f80b",
  1211 => x"80f52d71",
  1212 => x"82802905",
  1213 => x"80d7fa0b",
  1214 => x"80f52d70",
  1215 => x"84808029",
  1216 => x"1280d7fb",
  1217 => x"0b80f52d",
  1218 => x"7081800a",
  1219 => x"29127080",
  1220 => x"de8c0c80",
  1221 => x"de840871",
  1222 => x"2980ddf0",
  1223 => x"08057080",
  1224 => x"ddf40c80",
  1225 => x"d8810b80",
  1226 => x"f52d80d8",
  1227 => x"800b80f5",
  1228 => x"2d718280",
  1229 => x"290580d8",
  1230 => x"820b80f5",
  1231 => x"2d708480",
  1232 => x"80291280",
  1233 => x"d8830b80",
  1234 => x"f52d7098",
  1235 => x"2b81f00a",
  1236 => x"06720570",
  1237 => x"80ddf80c",
  1238 => x"80d8850b",
  1239 => x"80f52d80",
  1240 => x"d8840b80",
  1241 => x"f52d7188",
  1242 => x"2b075746",
  1243 => x"52575257",
  1244 => x"5d575152",
  1245 => x"5f525c57",
  1246 => x"57577580",
  1247 => x"de900b81",
  1248 => x"8a2dfe14",
  1249 => x"77297505",
  1250 => x"80ddfc0c",
  1251 => x"820b80d5",
  1252 => x"8c0c80dd",
  1253 => x"e008802e",
  1254 => x"81b93880",
  1255 => x"d7d45280",
  1256 => x"de940816",
  1257 => x"519cc22d",
  1258 => x"80d6f408",
  1259 => x"802e81a3",
  1260 => x"38845380",
  1261 => x"cfb85280",
  1262 => x"dbd0519e",
  1263 => x"e82d80d6",
  1264 => x"f408818f",
  1265 => x"3880dbbd",
  1266 => x"0b80f52d",
  1267 => x"80dbbc0b",
  1268 => x"80f52d71",
  1269 => x"882b0780",
  1270 => x"dbbe0b80",
  1271 => x"f52d7090",
  1272 => x"2b720780",
  1273 => x"dbbf0b80",
  1274 => x"f52d7098",
  1275 => x"2b720780",
  1276 => x"d58c0c5b",
  1277 => x"5258555a",
  1278 => x"a8d30480",
  1279 => x"d7e60b80",
  1280 => x"f52d80d7",
  1281 => x"e50b80f5",
  1282 => x"2d718280",
  1283 => x"29057080",
  1284 => x"dde40c70",
  1285 => x"a02983ff",
  1286 => x"0570892a",
  1287 => x"7080de80",
  1288 => x"0c80d7eb",
  1289 => x"0b80f52d",
  1290 => x"80d7ea0b",
  1291 => x"80f52d71",
  1292 => x"82802905",
  1293 => x"7080de8c",
  1294 => x"0c7b7129",
  1295 => x"1e7080dd",
  1296 => x"fc0c7d80",
  1297 => x"ddf80c73",
  1298 => x"0580ddf4",
  1299 => x"0c5a5451",
  1300 => x"51555980",
  1301 => x"519fde2d",
  1302 => x"81557480",
  1303 => x"d6f40c02",
  1304 => x"a8050d04",
  1305 => x"02f0050d",
  1306 => x"80d58808",
  1307 => x"53728025",
  1308 => x"80c73872",
  1309 => x"fe0a0653",
  1310 => x"72fe0a2e",
  1311 => x"b1388054",
  1312 => x"80de8408",
  1313 => x"742ea738",
  1314 => x"80dea452",
  1315 => x"80d58808",
  1316 => x"fe0a0680",
  1317 => x"ddf00805",
  1318 => x"7480de8c",
  1319 => x"08290551",
  1320 => x"9aff2d81",
  1321 => x"145480de",
  1322 => x"84087426",
  1323 => x"db3880d5",
  1324 => x"8808fe0a",
  1325 => x"0680d588",
  1326 => x"0c029005",
  1327 => x"0d0402f0",
  1328 => x"050d7570",
  1329 => x"872a5553",
  1330 => x"80dde008",
  1331 => x"85387288",
  1332 => x"2a5480d5",
  1333 => x"8808fe0a",
  1334 => x"06537373",
  1335 => x"2ea338a8",
  1336 => x"e42d80de",
  1337 => x"a45280dd",
  1338 => x"f0081451",
  1339 => x"9cc22d80",
  1340 => x"d6f40853",
  1341 => x"80d6f408",
  1342 => x"802e8838",
  1343 => x"7380d588",
  1344 => x"0c815372",
  1345 => x"80d6f40c",
  1346 => x"0290050d",
  1347 => x"0402f405",
  1348 => x"0d747052",
  1349 => x"53a9be2d",
  1350 => x"80d6f408",
  1351 => x"5280d6f4",
  1352 => x"08802e8b",
  1353 => x"3872519f",
  1354 => x"a72d80d6",
  1355 => x"f4085271",
  1356 => x"80d6f40c",
  1357 => x"028c050d",
  1358 => x"0402f805",
  1359 => x"0d735271",
  1360 => x"51a9be2d",
  1361 => x"80d6f408",
  1362 => x"893880d6",
  1363 => x"f40852aa",
  1364 => x"e5047151",
  1365 => x"9fa72d80",
  1366 => x"d6f40880",
  1367 => x"2e873881",
  1368 => x"1252aabf",
  1369 => x"047180d6",
  1370 => x"f40c0288",
  1371 => x"050d0402",
  1372 => x"f4050d74",
  1373 => x"80dde008",
  1374 => x"52537080",
  1375 => x"2e9e3880",
  1376 => x"7380ffff",
  1377 => x"fff80652",
  1378 => x"527080ff",
  1379 => x"fffff82e",
  1380 => x"09810683",
  1381 => x"38815271",
  1382 => x"51aba804",
  1383 => x"7283ffff",
  1384 => x"2e098106",
  1385 => x"83388151",
  1386 => x"7080d6f4",
  1387 => x"0c028c05",
  1388 => x"0d0402f4",
  1389 => x"050d7476",
  1390 => x"71535452",
  1391 => x"a9be2d80",
  1392 => x"d6f40880",
  1393 => x"2e80c638",
  1394 => x"80dde008",
  1395 => x"802e9b38",
  1396 => x"71822b83",
  1397 => x"fc0680de",
  1398 => x"a4117453",
  1399 => x"5152be8a",
  1400 => x"2d80d6f4",
  1401 => x"08720cac",
  1402 => x"82047110",
  1403 => x"83fe0680",
  1404 => x"dea41174",
  1405 => x"535152be",
  1406 => x"b52d80d6",
  1407 => x"f4087281",
  1408 => x"8a2d80d5",
  1409 => x"8808810a",
  1410 => x"0780d588",
  1411 => x"0c028c05",
  1412 => x"0d0402dc",
  1413 => x"050d7b80",
  1414 => x"ddd80884",
  1415 => x"80291cff",
  1416 => x"11892a70",
  1417 => x"80de8808",
  1418 => x"2a705a5a",
  1419 => x"515559fe",
  1420 => x"0a0b80d5",
  1421 => x"880c80d5",
  1422 => x"8c0851aa",
  1423 => x"b92d80d6",
  1424 => x"f40880d6",
  1425 => x"f4085955",
  1426 => x"817725a0",
  1427 => x"38811551",
  1428 => x"aab92d80",
  1429 => x"d6f40880",
  1430 => x"d6f40853",
  1431 => x"755254ab",
  1432 => x"b22d73ff",
  1433 => x"17575575",
  1434 => x"8124e238",
  1435 => x"f00a5480",
  1436 => x"dde00885",
  1437 => x"3883ffff",
  1438 => x"54735274",
  1439 => x"51abb22d",
  1440 => x"78802e88",
  1441 => x"38775278",
  1442 => x"51abb22d",
  1443 => x"a8e42d76",
  1444 => x"09810555",
  1445 => x"80dde008",
  1446 => x"802e81aa",
  1447 => x"3880d7d4",
  1448 => x"5280de90",
  1449 => x"0b80e02d",
  1450 => x"80de9408",
  1451 => x"05519cc2",
  1452 => x"2d80d6f4",
  1453 => x"08802e81",
  1454 => x"8d388453",
  1455 => x"80cfb852",
  1456 => x"80dbd051",
  1457 => x"9ee82d80",
  1458 => x"d6f40880",
  1459 => x"f93880db",
  1460 => x"bd0b80f5",
  1461 => x"2d80dbbc",
  1462 => x"0b80f52d",
  1463 => x"71882b07",
  1464 => x"80dbbe0b",
  1465 => x"80f52d70",
  1466 => x"902b7207",
  1467 => x"80dbbf0b",
  1468 => x"80f52d70",
  1469 => x"982b7207",
  1470 => x"7a115152",
  1471 => x"5b525255",
  1472 => x"567380db",
  1473 => x"bc0b81b7",
  1474 => x"2d73882a",
  1475 => x"557480db",
  1476 => x"bd0b81b7",
  1477 => x"2d73902a",
  1478 => x"557480db",
  1479 => x"be0b81b7",
  1480 => x"2d73982a",
  1481 => x"557480db",
  1482 => x"bf0b81b7",
  1483 => x"2d7380d5",
  1484 => x"8c0c80d7",
  1485 => x"d45280de",
  1486 => x"900b80e0",
  1487 => x"2d80de94",
  1488 => x"0805519a",
  1489 => x"ff2d7780",
  1490 => x"d6f40c02",
  1491 => x"a4050d04",
  1492 => x"02ec050d",
  1493 => x"76558070",
  1494 => x"7680f52d",
  1495 => x"53545270",
  1496 => x"722e8338",
  1497 => x"81537081",
  1498 => x"e52e9f38",
  1499 => x"81707406",
  1500 => x"52547080",
  1501 => x"2e94388b",
  1502 => x"1580f52d",
  1503 => x"70832a70",
  1504 => x"76065152",
  1505 => x"55708338",
  1506 => x"73527180",
  1507 => x"d6f40c02",
  1508 => x"94050d04",
  1509 => x"02e4050d",
  1510 => x"7970842c",
  1511 => x"1a718f06",
  1512 => x"52555372",
  1513 => x"8a3880d7",
  1514 => x"d4527351",
  1515 => x"9cc22d72",
  1516 => x"a02980d7",
  1517 => x"d4055480",
  1518 => x"7480f52d",
  1519 => x"56537473",
  1520 => x"2e833881",
  1521 => x"537481e5",
  1522 => x"2e81f138",
  1523 => x"72802e81",
  1524 => x"eb388b14",
  1525 => x"80f52d70",
  1526 => x"832a8106",
  1527 => x"58567699",
  1528 => x"3880d584",
  1529 => x"08537289",
  1530 => x"387280db",
  1531 => x"d40b81b7",
  1532 => x"2d7680d5",
  1533 => x"840cb1bc",
  1534 => x"04758f2e",
  1535 => x"09810681",
  1536 => x"bb38749f",
  1537 => x"068d2980",
  1538 => x"dbc71151",
  1539 => x"53811480",
  1540 => x"f52d7370",
  1541 => x"81055581",
  1542 => x"b72d8314",
  1543 => x"80f52d73",
  1544 => x"70810555",
  1545 => x"81b72d85",
  1546 => x"1480f52d",
  1547 => x"73708105",
  1548 => x"5581b72d",
  1549 => x"871480f5",
  1550 => x"2d737081",
  1551 => x"055581b7",
  1552 => x"2d891480",
  1553 => x"f52d7370",
  1554 => x"81055581",
  1555 => x"b72d8e14",
  1556 => x"80f52d73",
  1557 => x"70810555",
  1558 => x"81b72d90",
  1559 => x"1480f52d",
  1560 => x"73708105",
  1561 => x"5581b72d",
  1562 => x"921480f5",
  1563 => x"2d737081",
  1564 => x"055581b7",
  1565 => x"2d941480",
  1566 => x"f52d7370",
  1567 => x"81055581",
  1568 => x"b72d9614",
  1569 => x"80f52d73",
  1570 => x"70810555",
  1571 => x"81b72d98",
  1572 => x"1480f52d",
  1573 => x"73708105",
  1574 => x"5581b72d",
  1575 => x"9c1480f5",
  1576 => x"2d737081",
  1577 => x"055581b7",
  1578 => x"2d9e1480",
  1579 => x"f52d7381",
  1580 => x"b72d80d5",
  1581 => x"84088105",
  1582 => x"80d5840c",
  1583 => x"7380d6f4",
  1584 => x"0c029c05",
  1585 => x"0d0402e0",
  1586 => x"050d797b",
  1587 => x"59578070",
  1588 => x"5752b293",
  1589 => x"0473ae2e",
  1590 => x"09810694",
  1591 => x"38718724",
  1592 => x"af387612",
  1593 => x"51a07181",
  1594 => x"b72d8112",
  1595 => x"52b1dd04",
  1596 => x"76125572",
  1597 => x"8113ff9f",
  1598 => x"157081ff",
  1599 => x"06515353",
  1600 => x"54709926",
  1601 => x"86387281",
  1602 => x"df065473",
  1603 => x"7581b72d",
  1604 => x"81165680",
  1605 => x"76197080",
  1606 => x"f52d7081",
  1607 => x"ff065755",
  1608 => x"52557375",
  1609 => x"2e833881",
  1610 => x"55718a24",
  1611 => x"983874ff",
  1612 => x"a438718a",
  1613 => x"248f3876",
  1614 => x"1251a071",
  1615 => x"81b72d81",
  1616 => x"1252b2b2",
  1617 => x"04800b8b",
  1618 => x"1881b72d",
  1619 => x"02a0050d",
  1620 => x"0402ec05",
  1621 => x"0d76789c",
  1622 => x"11085355",
  1623 => x"55be8a2d",
  1624 => x"80d6f408",
  1625 => x"84160c9a",
  1626 => x"1480e02d",
  1627 => x"51beb52d",
  1628 => x"80d6f408",
  1629 => x"80d6f408",
  1630 => x"88170c80",
  1631 => x"d6f40853",
  1632 => x"5380dde0",
  1633 => x"08802e99",
  1634 => x"38941480",
  1635 => x"e02d51be",
  1636 => x"b52d80d6",
  1637 => x"f408902b",
  1638 => x"83fff00a",
  1639 => x"06701451",
  1640 => x"52718816",
  1641 => x"0c80750c",
  1642 => x"810b80d6",
  1643 => x"f40c0294",
  1644 => x"050d0402",
  1645 => x"d4050d7d",
  1646 => x"5b807080",
  1647 => x"de980856",
  1648 => x"575a7380",
  1649 => x"ddf8082e",
  1650 => x"09810683",
  1651 => x"38815a73",
  1652 => x"80de9c08",
  1653 => x"56578059",
  1654 => x"80dde408",
  1655 => x"792e80e9",
  1656 => x"38788f06",
  1657 => x"a0175754",
  1658 => x"73913880",
  1659 => x"d7d45274",
  1660 => x"51811555",
  1661 => x"9cc22d80",
  1662 => x"d7d45680",
  1663 => x"7680f52d",
  1664 => x"55587378",
  1665 => x"2e833881",
  1666 => x"587381e5",
  1667 => x"2eaf3877",
  1668 => x"802eaa38",
  1669 => x"8b1680f5",
  1670 => x"2d980654",
  1671 => x"739f388b",
  1672 => x"537a5275",
  1673 => x"519ee82d",
  1674 => x"80d6f408",
  1675 => x"90387552",
  1676 => x"7c51b2d1",
  1677 => x"2d80d6f4",
  1678 => x"0854b4f8",
  1679 => x"04811959",
  1680 => x"80dde408",
  1681 => x"7926ff99",
  1682 => x"3879802e",
  1683 => x"a9387651",
  1684 => x"aa8d2d80",
  1685 => x"d6f40880",
  1686 => x"d6f40852",
  1687 => x"57aaef2d",
  1688 => x"80d6f408",
  1689 => x"9138fe17",
  1690 => x"80ddd808",
  1691 => x"2980ddf4",
  1692 => x"080555b3",
  1693 => x"d6048054",
  1694 => x"7380d6f4",
  1695 => x"0c02ac05",
  1696 => x"0d0402f4",
  1697 => x"050d7470",
  1698 => x"08810571",
  1699 => x"0c700880",
  1700 => x"dddc0806",
  1701 => x"5353718f",
  1702 => x"38881308",
  1703 => x"51aa8d2d",
  1704 => x"80d6f408",
  1705 => x"88140c81",
  1706 => x"0b80d6f4",
  1707 => x"0c028c05",
  1708 => x"0d0402f0",
  1709 => x"050d7588",
  1710 => x"1108fe05",
  1711 => x"80ddd808",
  1712 => x"2980ddf4",
  1713 => x"08057108",
  1714 => x"80dddc08",
  1715 => x"060580d6",
  1716 => x"f40c5402",
  1717 => x"90050d04",
  1718 => x"02f0050d",
  1719 => x"75881108",
  1720 => x"fe0580dd",
  1721 => x"d8082980",
  1722 => x"ddf40811",
  1723 => x"720880dd",
  1724 => x"dc080605",
  1725 => x"79555354",
  1726 => x"549aff2d",
  1727 => x"0290050d",
  1728 => x"0402ffbc",
  1729 => x"050d6264",
  1730 => x"66686a43",
  1731 => x"43435a5a",
  1732 => x"80707172",
  1733 => x"415e5e5b",
  1734 => x"7980ddf8",
  1735 => x"082e0981",
  1736 => x"06893880",
  1737 => x"dde0087b",
  1738 => x"2e833881",
  1739 => x"5e805780",
  1740 => x"dde40877",
  1741 => x"2e819338",
  1742 => x"76527851",
  1743 => x"af942d80",
  1744 => x"d6f40856",
  1745 => x"7e913880",
  1746 => x"d6f40851",
  1747 => x"aed02d80",
  1748 => x"d6f40880",
  1749 => x"2ebb387c",
  1750 => x"55761b54",
  1751 => x"80dbd453",
  1752 => x"75526051",
  1753 => x"7f2d80d6",
  1754 => x"f4088025",
  1755 => x"8638815c",
  1756 => x"b7910480",
  1757 => x"0b80d6f4",
  1758 => x"08259638",
  1759 => x"7b802e80",
  1760 => x"c93880d7",
  1761 => x"d4527684",
  1762 => x"2c19519a",
  1763 => x"ff2db7ca",
  1764 => x"0480d584",
  1765 => x"085d8077",
  1766 => x"8f065758",
  1767 => x"758f2e09",
  1768 => x"81068338",
  1769 => x"81587b80",
  1770 => x"2e943877",
  1771 => x"802e8f38",
  1772 => x"80d7d452",
  1773 => x"76842c19",
  1774 => x"519aff2d",
  1775 => x"805c8117",
  1776 => x"5780dde4",
  1777 => x"087726fe",
  1778 => x"ef3880dd",
  1779 => x"e4087726",
  1780 => x"b4387d80",
  1781 => x"2eaf3879",
  1782 => x"51aa8d2d",
  1783 => x"80d6f408",
  1784 => x"80d6f408",
  1785 => x"525aaaef",
  1786 => x"2d80d6f4",
  1787 => x"089738fe",
  1788 => x"1a80ddd8",
  1789 => x"082980dd",
  1790 => x"f4080580",
  1791 => x"dde4081c",
  1792 => x"5c59b6ad",
  1793 => x"040280c4",
  1794 => x"050d0402",
  1795 => x"ec050d78",
  1796 => x"55775476",
  1797 => x"5380de9c",
  1798 => x"085280de",
  1799 => x"980851b6",
  1800 => x"812d0294",
  1801 => x"050d0402",
  1802 => x"e8050d77",
  1803 => x"797c5856",
  1804 => x"5474802e",
  1805 => x"bc388853",
  1806 => x"84145274",
  1807 => x"519ee82d",
  1808 => x"80d6f408",
  1809 => x"ac388353",
  1810 => x"8c145288",
  1811 => x"15519ee8",
  1812 => x"2d80d6f4",
  1813 => x"089b3881",
  1814 => x"740c7494",
  1815 => x"150c757c",
  1816 => x"3198150c",
  1817 => x"759c150c",
  1818 => x"7990150c",
  1819 => x"8154b8f3",
  1820 => x"04805473",
  1821 => x"80d6f40c",
  1822 => x"0298050d",
  1823 => x"0402c805",
  1824 => x"0d606053",
  1825 => x"02bc05e4",
  1826 => x"055256b1",
  1827 => x"c62d8057",
  1828 => x"8053b8a7",
  1829 => x"5202b805",
  1830 => x"e00551b8",
  1831 => x"8b2d7580",
  1832 => x"2ea6387b",
  1833 => x"941180e0",
  1834 => x"2d5254be",
  1835 => x"b52d80d6",
  1836 => x"f408902b",
  1837 => x"7c9a1180",
  1838 => x"e02d5355",
  1839 => x"55beb52d",
  1840 => x"7480d6f4",
  1841 => x"0807760c",
  1842 => x"7680d6f4",
  1843 => x"0c02b805",
  1844 => x"0d0402f8",
  1845 => x"050d8052",
  1846 => x"7351b8fd",
  1847 => x"2d028805",
  1848 => x"0d0402f8",
  1849 => x"050d8075",
  1850 => x"7080f52d",
  1851 => x"51525270",
  1852 => x"81e52e09",
  1853 => x"81068338",
  1854 => x"81527009",
  1855 => x"81057080",
  1856 => x"25730770",
  1857 => x"54515170",
  1858 => x"802e8838",
  1859 => x"7377710c",
  1860 => x"51815271",
  1861 => x"80d6f40c",
  1862 => x"0288050d",
  1863 => x"0402e005",
  1864 => x"0d797b9c",
  1865 => x"12085758",
  1866 => x"58815674",
  1867 => x"81aa3874",
  1868 => x"7780f52d",
  1869 => x"55567381",
  1870 => x"e52e0981",
  1871 => x"06833881",
  1872 => x"56730981",
  1873 => x"05708025",
  1874 => x"77077058",
  1875 => x"51547380",
  1876 => x"2e818538",
  1877 => x"88538418",
  1878 => x"52765180",
  1879 => x"ccfe2d83",
  1880 => x"538c1852",
  1881 => x"88175180",
  1882 => x"ccfe2d98",
  1883 => x"1880f52d",
  1884 => x"8b1881b7",
  1885 => x"2d748c18",
  1886 => x"81b72d74",
  1887 => x"8d1881b7",
  1888 => x"2d749618",
  1889 => x"818a2d74",
  1890 => x"8e18818a",
  1891 => x"2d749818",
  1892 => x"818a2d74",
  1893 => x"9018818a",
  1894 => x"2d749218",
  1895 => x"818a2d96",
  1896 => x"1880e02d",
  1897 => x"51beb52d",
  1898 => x"80d6f408",
  1899 => x"9a18818a",
  1900 => x"2d941880",
  1901 => x"e02d51be",
  1902 => x"b52d80d6",
  1903 => x"f4089418",
  1904 => x"818a2d90",
  1905 => x"180851be",
  1906 => x"8a2d80d6",
  1907 => x"f4089c18",
  1908 => x"0c810b9c",
  1909 => x"190cff56",
  1910 => x"7580d6f4",
  1911 => x"0c02a005",
  1912 => x"0d0402c0",
  1913 => x"050d6163",
  1914 => x"71535957",
  1915 => x"b9d22d80",
  1916 => x"5480d6f4",
  1917 => x"08742e09",
  1918 => x"810681e6",
  1919 => x"38bc8804",
  1920 => x"80d6f408",
  1921 => x"54bcd904",
  1922 => x"ff598153",
  1923 => x"b9e25202",
  1924 => x"a0057052",
  1925 => x"56b88b2d",
  1926 => x"78802581",
  1927 => x"8a3880dd",
  1928 => x"e008802e",
  1929 => x"81813880",
  1930 => x"de980854",
  1931 => x"7351a9be",
  1932 => x"2d80d6f4",
  1933 => x"08802ec8",
  1934 => x"3873519f",
  1935 => x"a72d80d6",
  1936 => x"f40851aa",
  1937 => x"ef2d80d6",
  1938 => x"f4088e38",
  1939 => x"73519fa7",
  1940 => x"2d80d6f4",
  1941 => x"0854bcac",
  1942 => x"04735281",
  1943 => x"51ac922d",
  1944 => x"80d6f408",
  1945 => x"fe0580dd",
  1946 => x"d8082980",
  1947 => x"ddf40805",
  1948 => x"55848053",
  1949 => x"805280d7",
  1950 => x"d45180cd",
  1951 => x"a92d8054",
  1952 => x"80ddd808",
  1953 => x"742e9638",
  1954 => x"80d7d452",
  1955 => x"7315519a",
  1956 => x"ff2d8114",
  1957 => x"5480ddd8",
  1958 => x"087426ec",
  1959 => x"388153b9",
  1960 => x"e2527551",
  1961 => x"b88b2d80",
  1962 => x"54737924",
  1963 => x"b5387652",
  1964 => x"0280c005",
  1965 => x"e40551b1",
  1966 => x"c62d775d",
  1967 => x"80527751",
  1968 => x"ac922d80",
  1969 => x"d6f4085e",
  1970 => x"8040a002",
  1971 => x"bc0581b7",
  1972 => x"2d8153ba",
  1973 => x"9d520280",
  1974 => x"c005e005",
  1975 => x"51b88b2d",
  1976 => x"7f547380",
  1977 => x"d6f40c02",
  1978 => x"80c0050d",
  1979 => x"0402f405",
  1980 => x"0d80de8c",
  1981 => x"0880ddd8",
  1982 => x"0829872b",
  1983 => x"80ddfc08",
  1984 => x"0580d6f4",
  1985 => x"0c028c05",
  1986 => x"0d0402f4",
  1987 => x"050d7470",
  1988 => x"882a83fe",
  1989 => x"80067072",
  1990 => x"982a0772",
  1991 => x"882b87fc",
  1992 => x"80800671",
  1993 => x"0773982b",
  1994 => x"0780d6f4",
  1995 => x"0c515351",
  1996 => x"028c050d",
  1997 => x"0402f805",
  1998 => x"0d028e05",
  1999 => x"80f52d74",
  2000 => x"882b0770",
  2001 => x"83ffff06",
  2002 => x"80d6f40c",
  2003 => x"51028805",
  2004 => x"0d0402f4",
  2005 => x"050d7476",
  2006 => x"78535452",
  2007 => x"80712597",
  2008 => x"38727081",
  2009 => x"055480f5",
  2010 => x"2d727081",
  2011 => x"055481b7",
  2012 => x"2dff1151",
  2013 => x"70eb3880",
  2014 => x"7281b72d",
  2015 => x"028c050d",
  2016 => x"0402dc05",
  2017 => x"0d7a7c71",
  2018 => x"08565a56",
  2019 => x"73802e89",
  2020 => x"38ff1476",
  2021 => x"0c80c0ed",
  2022 => x"04841608",
  2023 => x"55815474",
  2024 => x"8b2481cb",
  2025 => x"388b1980",
  2026 => x"f52d7084",
  2027 => x"2a708106",
  2028 => x"771080db",
  2029 => x"d40b80f5",
  2030 => x"2d5c5351",
  2031 => x"55577380",
  2032 => x"2e80e838",
  2033 => x"7417822b",
  2034 => x"80c39b0b",
  2035 => x"80d59812",
  2036 => x"0c548416",
  2037 => x"08902984",
  2038 => x"17083170",
  2039 => x"1080e2a8",
  2040 => x"05515490",
  2041 => x"7481b72d",
  2042 => x"84160890",
  2043 => x"29841708",
  2044 => x"31701080",
  2045 => x"e2a90551",
  2046 => x"54a07481",
  2047 => x"b72d7781",
  2048 => x"ff068417",
  2049 => x"08565473",
  2050 => x"802e8b38",
  2051 => x"9c5380db",
  2052 => x"d45280c0",
  2053 => x"9a048b53",
  2054 => x"78527490",
  2055 => x"29753170",
  2056 => x"1080e2aa",
  2057 => x"05525480",
  2058 => x"c0e20474",
  2059 => x"17822b80",
  2060 => x"c19a0b80",
  2061 => x"d598120c",
  2062 => x"547781ff",
  2063 => x"06841708",
  2064 => x"56547380",
  2065 => x"2e8b389c",
  2066 => x"5380dbd4",
  2067 => x"5280c0d5",
  2068 => x"048b5378",
  2069 => x"52749029",
  2070 => x"75317010",
  2071 => x"80e2a805",
  2072 => x"52548416",
  2073 => x"08810584",
  2074 => x"170cbed2",
  2075 => x"2d805473",
  2076 => x"80d6f40c",
  2077 => x"02a4050d",
  2078 => x"0402e805",
  2079 => x"0d775580",
  2080 => x"56805380",
  2081 => x"c3cb5202",
  2082 => x"9805f805",
  2083 => x"51b88b2d",
  2084 => x"7580d6f4",
  2085 => x"0c029805",
  2086 => x"0d0402ec",
  2087 => x"050d80d6",
  2088 => x"c4081751",
  2089 => x"80c0f92d",
  2090 => x"80d6f408",
  2091 => x"5580d6f4",
  2092 => x"08802ea1",
  2093 => x"388b5380",
  2094 => x"d6f40852",
  2095 => x"80dbd451",
  2096 => x"bed22d80",
  2097 => x"e2a40854",
  2098 => x"73802e89",
  2099 => x"38745280",
  2100 => x"dbd45173",
  2101 => x"2d029405",
  2102 => x"0d0402e0",
  2103 => x"050d80d6",
  2104 => x"c4085780",
  2105 => x"588053bf",
  2106 => x"815202a0",
  2107 => x"05f80551",
  2108 => x"b88b2d77",
  2109 => x"55748b24",
  2110 => x"a2387490",
  2111 => x"29753170",
  2112 => x"1080e2a8",
  2113 => x"05575480",
  2114 => x"7681b72d",
  2115 => x"9e168116",
  2116 => x"70575556",
  2117 => x"8b7425ef",
  2118 => x"38735802",
  2119 => x"a0050d04",
  2120 => x"02fc050d",
  2121 => x"725170fd",
  2122 => x"2eb23870",
  2123 => x"fd248b38",
  2124 => x"70fc2e80",
  2125 => x"d03880c3",
  2126 => x"8f0470fe",
  2127 => x"2eb93870",
  2128 => x"ff2e0981",
  2129 => x"0680c838",
  2130 => x"80d6c408",
  2131 => x"5170802e",
  2132 => x"be38ff11",
  2133 => x"80d6c40c",
  2134 => x"80c38f04",
  2135 => x"80d6c408",
  2136 => x"f4057080",
  2137 => x"d6c40c51",
  2138 => x"708025a3",
  2139 => x"38800b80",
  2140 => x"d6c40c80",
  2141 => x"c38f0480",
  2142 => x"d6c40881",
  2143 => x"0580d6c4",
  2144 => x"0c80c38f",
  2145 => x"0480d6c4",
  2146 => x"088c0580",
  2147 => x"d6c40c80",
  2148 => x"c1da2d8f",
  2149 => x"df2d0284",
  2150 => x"050d0402",
  2151 => x"fc050d80",
  2152 => x"d6c40813",
  2153 => x"5180c0f9",
  2154 => x"2d80d6f4",
  2155 => x"08802e89",
  2156 => x"3880d6f4",
  2157 => x"08519fde",
  2158 => x"2d800b80",
  2159 => x"d6c40c80",
  2160 => x"c1da2d8f",
  2161 => x"df2d0284",
  2162 => x"050d0402",
  2163 => x"f4050d74",
  2164 => x"52807208",
  2165 => x"52537073",
  2166 => x"2e8938ff",
  2167 => x"11720c80",
  2168 => x"c3e90475",
  2169 => x"84130c81",
  2170 => x"537280d6",
  2171 => x"f40c028c",
  2172 => x"050d0402",
  2173 => x"fc050d80",
  2174 => x"0b80d6c4",
  2175 => x"0c80c1da",
  2176 => x"2d8fa02d",
  2177 => x"80d6f408",
  2178 => x"80d6b40c",
  2179 => x"80d59051",
  2180 => x"90cd2d02",
  2181 => x"84050d04",
  2182 => x"7180e2a4",
  2183 => x"0c0402f8",
  2184 => x"050dff14",
  2185 => x"51805270",
  2186 => x"722e8b38",
  2187 => x"81127181",
  2188 => x"2c525270",
  2189 => x"f738f712",
  2190 => x"80d6f40c",
  2191 => x"0288050d",
  2192 => x"0402c405",
  2193 => x"0d606264",
  2194 => x"72545659",
  2195 => x"55b9d22d",
  2196 => x"805380d6",
  2197 => x"f408732e",
  2198 => x"09810681",
  2199 => x"8c387352",
  2200 => x"7451bbe2",
  2201 => x"2d80d6f4",
  2202 => x"085380d6",
  2203 => x"f408802e",
  2204 => x"80f73881",
  2205 => x"5377802e",
  2206 => x"80ef3880",
  2207 => x"74525680",
  2208 => x"c49e2d80",
  2209 => x"d6f40875",
  2210 => x"5302a405",
  2211 => x"70535457",
  2212 => x"b1c62d72",
  2213 => x"5202bc05",
  2214 => x"f40551b3",
  2215 => x"b32d80d6",
  2216 => x"f4085380",
  2217 => x"d6f40876",
  2218 => x"2ebf3875",
  2219 => x"7425b838",
  2220 => x"76527551",
  2221 => x"84c32d80",
  2222 => x"d7d45177",
  2223 => x"2d80d6f4",
  2224 => x"08802e8e",
  2225 => x"3880d7d4",
  2226 => x"5202bc05",
  2227 => x"f40551b5",
  2228 => x"d82d02bc",
  2229 => x"05f40551",
  2230 => x"b5822dfc",
  2231 => x"80148117",
  2232 => x"57547380",
  2233 => x"24ca3881",
  2234 => x"537280d6",
  2235 => x"f40c02bc",
  2236 => x"050d0402",
  2237 => x"c8050d60",
  2238 => x"6202b405",
  2239 => x"56585372",
  2240 => x"802e8c38",
  2241 => x"72527351",
  2242 => x"b2d12d80",
  2243 => x"c6a1047f",
  2244 => x"52029c05",
  2245 => x"705253b1",
  2246 => x"c62d7252",
  2247 => x"7351b3b3",
  2248 => x"2d80d6f4",
  2249 => x"085480d6",
  2250 => x"f408802e",
  2251 => x"bf387c54",
  2252 => x"80745255",
  2253 => x"80c49e2d",
  2254 => x"80d6f408",
  2255 => x"56747425",
  2256 => x"a9387552",
  2257 => x"745184c3",
  2258 => x"2d02ac05",
  2259 => x"705253b5",
  2260 => x"b22d80d6",
  2261 => x"f4085176",
  2262 => x"2d7251b5",
  2263 => x"822dfc80",
  2264 => x"14811656",
  2265 => x"54738024",
  2266 => x"d9387c54",
  2267 => x"7380d6f4",
  2268 => x"0c02b805",
  2269 => x"0d0402f0",
  2270 => x"050d7570",
  2271 => x"9f06718c",
  2272 => x"2a7280d6",
  2273 => x"cc0c7284",
  2274 => x"2a81fe06",
  2275 => x"71810605",
  2276 => x"70832b71",
  2277 => x"1114ff11",
  2278 => x"51555751",
  2279 => x"54555180",
  2280 => x"d6c8088a",
  2281 => x"38711013",
  2282 => x"7411ff05",
  2283 => x"51517080",
  2284 => x"d6f40c02",
  2285 => x"90050d04",
  2286 => x"02f4050d",
  2287 => x"f4900870",
  2288 => x"80c88080",
  2289 => x"06535371",
  2290 => x"802eb438",
  2291 => x"7283ffff",
  2292 => x"065180c6",
  2293 => x"f62d80d6",
  2294 => x"f40880d6",
  2295 => x"e80c800b",
  2296 => x"80d6dc0b",
  2297 => x"818a2d72",
  2298 => x"942a7081",
  2299 => x"06515271",
  2300 => x"802e8c38",
  2301 => x"80d6f408",
  2302 => x"810a0780",
  2303 => x"d6e80c72",
  2304 => x"81908080",
  2305 => x"06527180",
  2306 => x"2eb43872",
  2307 => x"83ffff06",
  2308 => x"5180c6f6",
  2309 => x"2d80d6f4",
  2310 => x"0880d6ec",
  2311 => x"0c800b80",
  2312 => x"d6de0b81",
  2313 => x"8a2d7295",
  2314 => x"2a708106",
  2315 => x"51527180",
  2316 => x"2e8c3880",
  2317 => x"d6f40881",
  2318 => x"0a0780d6",
  2319 => x"ec0c7290",
  2320 => x"2a708106",
  2321 => x"51527180",
  2322 => x"2e8f3880",
  2323 => x"d6d008e7",
  2324 => x"067080d6",
  2325 => x"d00cf490",
  2326 => x"0c028c05",
  2327 => x"0d0402e4",
  2328 => x"050d7870",
  2329 => x"822b80d6",
  2330 => x"e8117008",
  2331 => x"57575856",
  2332 => x"73ff2e81",
  2333 => x"e23873fe",
  2334 => x"0a06538c",
  2335 => x"c0732792",
  2336 => x"38ff750c",
  2337 => x"80d6d008",
  2338 => x"980780d6",
  2339 => x"d00c80ca",
  2340 => x"d704758c",
  2341 => x"c0291470",
  2342 => x"842980e5",
  2343 => x"b0057008",
  2344 => x"565153bd",
  2345 => x"ed2d7380",
  2346 => x"d6f40827",
  2347 => x"81983880",
  2348 => x"d7d45273",
  2349 => x"519cc22d",
  2350 => x"80d6f408",
  2351 => x"802e8186",
  2352 => x"38740880",
  2353 => x"2580c138",
  2354 => x"751080d6",
  2355 => x"dc057080",
  2356 => x"e02d80d7",
  2357 => x"d4055753",
  2358 => x"83ff55f4",
  2359 => x"94085372",
  2360 => x"76708105",
  2361 => x"5881b72d",
  2362 => x"84800bf4",
  2363 => x"940c800b",
  2364 => x"f4940cff",
  2365 => x"15557480",
  2366 => x"25e13880",
  2367 => x"d7d45273",
  2368 => x"519aff2d",
  2369 => x"80cab804",
  2370 => x"751080d6",
  2371 => x"dc057080",
  2372 => x"e02d80d7",
  2373 => x"d4055553",
  2374 => x"83ff5573",
  2375 => x"80f52d82",
  2376 => x"8007f494",
  2377 => x"0c737081",
  2378 => x"055580f5",
  2379 => x"2df4940c",
  2380 => x"ff155574",
  2381 => x"8025e438",
  2382 => x"80d6d008",
  2383 => x"900780d6",
  2384 => x"d00c80ca",
  2385 => x"d00480d6",
  2386 => x"d0089807",
  2387 => x"80d6d00c",
  2388 => x"ff0b80d6",
  2389 => x"e8180c02",
  2390 => x"9c050d04",
  2391 => x"02fc050d",
  2392 => x"80c7b82d",
  2393 => x"805180c8",
  2394 => x"de2d8151",
  2395 => x"80c8de2d",
  2396 => x"80d6d008",
  2397 => x"f4900c02",
  2398 => x"84050d04",
  2399 => x"02f4050d",
  2400 => x"80d6d408",
  2401 => x"8cc02980",
  2402 => x"d6d80805",
  2403 => x"70842980",
  2404 => x"e5b00576",
  2405 => x"710c5153",
  2406 => x"80d6d808",
  2407 => x"810580d6",
  2408 => x"d80c028c",
  2409 => x"050d0402",
  2410 => x"ec050d76",
  2411 => x"7080d6d4",
  2412 => x"0c55800b",
  2413 => x"80d6d80c",
  2414 => x"80cafc53",
  2415 => x"78527751",
  2416 => x"80c5f32d",
  2417 => x"80d6f408",
  2418 => x"09810570",
  2419 => x"80d6f408",
  2420 => x"079f2a51",
  2421 => x"547380d6",
  2422 => x"f01681b7",
  2423 => x"2d80d6f4",
  2424 => x"08ad8080",
  2425 => x"32700981",
  2426 => x"05707207",
  2427 => x"802580d6",
  2428 => x"c80c5555",
  2429 => x"80d6f408",
  2430 => x"5480d6f4",
  2431 => x"08802e83",
  2432 => x"38815473",
  2433 => x"80d6f40c",
  2434 => x"0294050d",
  2435 => x"0402e405",
  2436 => x"0d800b80",
  2437 => x"d6dc7158",
  2438 => x"5855800b",
  2439 => x"80d6f016",
  2440 => x"81b72d74",
  2441 => x"822b53ff",
  2442 => x"0b80d6e8",
  2443 => x"140cff0b",
  2444 => x"80d6e014",
  2445 => x"0c807781",
  2446 => x"8a2d80e5",
  2447 => x"b016548c",
  2448 => x"bf538074",
  2449 => x"70840556",
  2450 => x"0cff1353",
  2451 => x"728025f2",
  2452 => x"388115b2",
  2453 => x"80178219",
  2454 => x"59575581",
  2455 => x"7525ffba",
  2456 => x"38800b80",
  2457 => x"d6d80c80",
  2458 => x"0b80d6d4",
  2459 => x"0c800b80",
  2460 => x"d6d00c80",
  2461 => x"0b80d6cc",
  2462 => x"0c029c05",
  2463 => x"0d0402e8",
  2464 => x"050d7779",
  2465 => x"7b565656",
  2466 => x"80537274",
  2467 => x"25963872",
  2468 => x"16731652",
  2469 => x"527080f5",
  2470 => x"2d7281b7",
  2471 => x"2d811353",
  2472 => x"80cd8a04",
  2473 => x"0298050d",
  2474 => x"0402ec05",
  2475 => x"0d767902",
  2476 => x"88059f05",
  2477 => x"80f52d55",
  2478 => x"55558052",
  2479 => x"71742590",
  2480 => x"38711551",
  2481 => x"727181b7",
  2482 => x"2d811252",
  2483 => x"80cdbc04",
  2484 => x"0294050d",
  2485 => x"0402f405",
  2486 => x"0d747653",
  2487 => x"53717081",
  2488 => x"055380f5",
  2489 => x"2d517073",
  2490 => x"70810555",
  2491 => x"81b72d70",
  2492 => x"ec38028c",
  2493 => x"050d0402",
  2494 => x"f4050d74",
  2495 => x"76545271",
  2496 => x"70810553",
  2497 => x"80f52d51",
  2498 => x"70f538ff",
  2499 => x"12527270",
  2500 => x"81055480",
  2501 => x"f52d5170",
  2502 => x"72708105",
  2503 => x"5481b72d",
  2504 => x"70ec3802",
  2505 => x"8c050d04",
  2506 => x"02d0050d",
  2507 => x"7d7f5859",
  2508 => x"885380df",
  2509 => x"5202a405",
  2510 => x"70525880",
  2511 => x"cda92d80",
  2512 => x"02b00581",
  2513 => x"b72d8756",
  2514 => x"7518778f",
  2515 => x"06555580",
  2516 => x"d2cc1480",
  2517 => x"f52d7581",
  2518 => x"b72d7684",
  2519 => x"2cff1757",
  2520 => x"57758424",
  2521 => x"e3388079",
  2522 => x"80f52d55",
  2523 => x"5673762e",
  2524 => x"a2387518",
  2525 => x"761a5555",
  2526 => x"7380f52d",
  2527 => x"7581b72d",
  2528 => x"81165675",
  2529 => x"84248c38",
  2530 => x"75197080",
  2531 => x"f52d5154",
  2532 => x"73e03889",
  2533 => x"5302b005",
  2534 => x"f4055278",
  2535 => x"5180ccfe",
  2536 => x"2d02b005",
  2537 => x"0d040000",
  2538 => x"00ffffff",
  2539 => x"ff00ffff",
  2540 => x"ffff00ff",
  2541 => x"ffffff00",
  2542 => x"000055aa",
  2543 => x"00000000",
  2544 => x"496e7365",
  2545 => x"72742064",
  2546 => x"69736b20",
  2547 => x"30000000",
  2548 => x"57726974",
  2549 => x"65207072",
  2550 => x"6f746563",
  2551 => x"74206469",
  2552 => x"736b2030",
  2553 => x"00000000",
  2554 => x"496e7365",
  2555 => x"72742064",
  2556 => x"69736b20",
  2557 => x"31000000",
  2558 => x"57726974",
  2559 => x"65207072",
  2560 => x"6f746563",
  2561 => x"74206469",
  2562 => x"736b2031",
  2563 => x"00000000",
  2564 => x"43726561",
  2565 => x"74652062",
  2566 => x"6c616e6b",
  2567 => x"20646973",
  2568 => x"6b000000",
  2569 => x"4261636b",
  2570 => x"00000000",
  2571 => x"4469736b",
  2572 => x"206d656e",
  2573 => x"75202020",
  2574 => x"20202020",
  2575 => x"20202020",
  2576 => x"20100000",
  2577 => x"45786974",
  2578 => x"00000000",
  2579 => x"4469736b",
  2580 => x"206d656e",
  2581 => x"752e0000",
  2582 => x"4c6f6164",
  2583 => x"696e6720",
  2584 => x"6661696c",
  2585 => x"65640000",
  2586 => x"4f4b0000",
  2587 => x"4449534b",
  2588 => x"00000000",
  2589 => x"2e44534b",
  2590 => x"00000000",
  2591 => x"43726561",
  2592 => x"74696e67",
  2593 => x"2066696c",
  2594 => x"653a2000",
  2595 => x"496e6974",
  2596 => x"69616c69",
  2597 => x"7a696e67",
  2598 => x"20534420",
  2599 => x"63617264",
  2600 => x"0a000000",
  2601 => x"14200000",
  2602 => x"15200000",
  2603 => x"53442069",
  2604 => x"6e69742e",
  2605 => x"2e2e0a00",
  2606 => x"53442063",
  2607 => x"61726420",
  2608 => x"72657365",
  2609 => x"74206661",
  2610 => x"696c6564",
  2611 => x"210a0000",
  2612 => x"53444843",
  2613 => x"20657272",
  2614 => x"6f72210a",
  2615 => x"00000000",
  2616 => x"57726974",
  2617 => x"65206661",
  2618 => x"696c6564",
  2619 => x"0a000000",
  2620 => x"52656164",
  2621 => x"20666169",
  2622 => x"6c65640a",
  2623 => x"00000000",
  2624 => x"43617264",
  2625 => x"20696e69",
  2626 => x"74206661",
  2627 => x"696c6564",
  2628 => x"0a000000",
  2629 => x"46415431",
  2630 => x"36202020",
  2631 => x"00000000",
  2632 => x"46415433",
  2633 => x"32202020",
  2634 => x"00000000",
  2635 => x"4e6f2070",
  2636 => x"61727469",
  2637 => x"74696f6e",
  2638 => x"20736967",
  2639 => x"0a000000",
  2640 => x"42616420",
  2641 => x"70617274",
  2642 => x"0a000000",
  2643 => x"30313233",
  2644 => x"34353637",
  2645 => x"38396162",
  2646 => x"63646566",
  2647 => x"00000000",
  2648 => x"00000002",
  2649 => x"00000004",
  2650 => x"0000282c",
  2651 => x"00002988",
  2652 => x"00000002",
  2653 => x"00002844",
  2654 => x"000007a9",
  2655 => x"00000000",
  2656 => x"00000000",
  2657 => x"00000000",
  2658 => x"00000004",
  2659 => x"0000284c",
  2660 => x"00002988",
  2661 => x"00000004",
  2662 => x"000028dc",
  2663 => x"00002988",
  2664 => x"00000002",
  2665 => x"000027c0",
  2666 => x"00000379",
  2667 => x"00000001",
  2668 => x"000027d0",
  2669 => x"00000006",
  2670 => x"00000002",
  2671 => x"000027e8",
  2672 => x"00000398",
  2673 => x"00000001",
  2674 => x"000027f8",
  2675 => x"00000007",
  2676 => x"00000002",
  2677 => x"00002810",
  2678 => x"000003f0",
  2679 => x"00000004",
  2680 => x"000028dc",
  2681 => x"00002988",
  2682 => x"00000004",
  2683 => x"00002824",
  2684 => x"00002964",
  2685 => x"00000000",
  2686 => x"00000000",
  2687 => x"00000000",
  2688 => x"00000000",
  2689 => x"00000004",
  2690 => x"00002858",
  2691 => x"00002a04",
  2692 => x"00000004",
  2693 => x"00002868",
  2694 => x"00002964",
  2695 => x"00000000",
  2696 => x"00000000",
  2697 => x"00000000",
  2698 => x"00000000",
  2699 => x"00000000",
  2700 => x"00000000",
  2701 => x"00000000",
  2702 => x"00000000",
  2703 => x"00000000",
  2704 => x"00000000",
  2705 => x"00000000",
  2706 => x"00000000",
  2707 => x"00000000",
  2708 => x"00000000",
  2709 => x"00000000",
  2710 => x"00000000",
  2711 => x"00000000",
  2712 => x"00000000",
  2713 => x"00000000",
  2714 => x"00000000",
  2715 => x"00000000",
  2716 => x"00000000",
  2717 => x"00000000",
  2718 => x"00000000",
  2719 => x"000000c6",
  2720 => x"00000000",
  2721 => x"00000000",
  2722 => x"7fffffff",
  2723 => x"00000002",
  2724 => x"00000002",
  2725 => x"00003128",
  2726 => x"0000209a",
  2727 => x"00000002",
  2728 => x"00003146",
  2729 => x"0000209a",
  2730 => x"00000002",
  2731 => x"00003164",
  2732 => x"0000209a",
  2733 => x"00000002",
  2734 => x"00003182",
  2735 => x"0000209a",
  2736 => x"00000002",
  2737 => x"000031a0",
  2738 => x"0000209a",
  2739 => x"00000002",
  2740 => x"000031be",
  2741 => x"0000209a",
  2742 => x"00000002",
  2743 => x"000031dc",
  2744 => x"0000209a",
  2745 => x"00000002",
  2746 => x"000031fa",
  2747 => x"0000209a",
  2748 => x"00000002",
  2749 => x"00003218",
  2750 => x"0000209a",
  2751 => x"00000002",
  2752 => x"00003236",
  2753 => x"0000209a",
  2754 => x"00000002",
  2755 => x"00003254",
  2756 => x"0000209a",
  2757 => x"00000002",
  2758 => x"00003272",
  2759 => x"0000209a",
  2760 => x"00000002",
  2761 => x"00003290",
  2762 => x"0000209a",
  2763 => x"00000004",
  2764 => x"00002824",
  2765 => x"00000000",
  2766 => x"00000000",
  2767 => x"00000000",
  2768 => x"00002120",
  2769 => x"00000000",
  2770 => x"00000000",
  2771 => x"00000000",
  2772 => x"00000000",
  2773 => x"00000000",
  2774 => x"00000000",
  2775 => x"00000000",
  2776 => x"ffffffff",
  2777 => x"ffffffff",
  2778 => x"ffffffff",
  2779 => x"ffffffff",
  2780 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

