module keymap(input wire[13:0] addr, output reg[7:0] data);

always @* begin
  case(addr[13:0])
    16'h0035: data = 8'h03;
    16'h0036: data = 8'h40;
    16'h0038: data = 8'h70;
    16'h0039: data = 8'h27;
    16'h003A: data = 8'h80;
    16'h0046: data = 8'h01;
    16'h0047: data = 8'h10;
    16'h004B: data = 8'h04;
    16'h0051: data = 8'h08;
    16'h0052: data = 8'h01;
    16'h0053: data = 8'h08;
    16'h0055: data = 8'h02;
    16'h0056: data = 8'h01;
    16'h0059: data = 8'h03;
    16'h005A: data = 8'h01;
    16'h006A: data = 8'h02;
    16'h006D: data = 8'h01;
    16'h006E: data = 8'h02;
    16'h0071: data = 8'h01;
    16'h0072: data = 8'h01;
    16'h0075: data = 8'h02;
    16'h0076: data = 8'h02;
    16'h0079: data = 8'h03;
    16'h007A: data = 8'h02;
    16'h0086: data = 8'h08;
    16'h008A: data = 8'h04;
    16'h008D: data = 8'h01;
    16'h008E: data = 8'h04;
    16'h0091: data = 8'h02;
    16'h0092: data = 8'h04;
    16'h0095: data = 8'h03;
    16'h0096: data = 8'h08;
    16'h0099: data = 8'h03;
    16'h009A: data = 8'h04;
    16'h00A5: data = 8'h07;
    16'h00A6: data = 8'h01;
    16'h00AA: data = 8'h10;
    16'h00AD: data = 8'h01;
    16'h00AE: data = 8'h08;
    16'h00B1: data = 8'h02;
    16'h00B2: data = 8'h10;
    16'h00B5: data = 8'h02;
    16'h00B6: data = 8'h08;
    16'h00B9: data = 8'h03;
    16'h00BA: data = 8'h10;
    16'h00C5: data = 8'h07;
    16'h00C6: data = 8'h08;
    16'h00C9: data = 8'h07;
    16'h00CA: data = 8'h10;
    16'h00CD: data = 8'h06;
    16'h00CE: data = 8'h10;
    16'h00D1: data = 8'h01;
    16'h00D2: data = 8'h10;
    16'h00D5: data = 8'h05;
    16'h00D6: data = 8'h10;
    16'h00D9: data = 8'h04;
    16'h00DA: data = 8'h10;
    16'h00E9: data = 8'h07;
    16'h00EA: data = 8'h04;
    16'h00ED: data = 8'h06;
    16'h00EE: data = 8'h08;
    16'h00F1: data = 8'h05;
    16'h00F2: data = 8'h08;
    16'h00F5: data = 8'h04;
    16'h00F6: data = 8'h08;
    16'h00F9: data = 8'h04;
    16'h00FA: data = 8'h04;
    16'h0105: data = 8'h07;
    16'h0106: data = 8'h20;
    16'h0109: data = 8'h06;
    16'h010A: data = 8'h04;
    16'h010D: data = 8'h05;
    16'h010E: data = 8'h04;
    16'h0111: data = 8'h05;
    16'h0112: data = 8'h02;
    16'h0115: data = 8'h04;
    16'h0116: data = 8'h01;
    16'h0119: data = 8'h04;
    16'h011A: data = 8'h02;
    16'h0125: data = 8'h07;
    16'h0126: data = 8'h40;
    16'h0129: data = 8'h04;
    16'h012A: data = 8'h20;
    16'h012D: data = 8'h06;
    16'h012E: data = 8'h02;
    16'h0131: data = 8'h14;
    16'h0132: data = 8'h01;
    16'h0135: data = 8'h05;
    16'h0136: data = 8'h01;
    16'h0139: data = 8'h14;
    16'h013A: data = 8'h08;
    16'h0148: data = 8'h70;
    16'h0149: data = 8'h21;
    16'h014A: data = 8'h08;
    16'h0150: data = 8'h70;
    16'h0151: data = 8'h26;
    16'h0152: data = 8'h02;
    16'h0161: data = 8'h03;
    16'h0162: data = 8'h80;
    16'h0167: data = 8'h04;
    16'h0169: data = 8'h06;
    16'h016A: data = 8'h01;
    16'h016D: data = 8'h04;
    16'h016E: data = 8'h40;
    16'h0174: data = 8'h70;
    16'h0175: data = 8'h21;
    16'h0176: data = 8'h10;
    16'h0184: data = 8'h70;
    16'h0185: data = 8'h22;
    16'h0186: data = 8'h01;
    16'h0199: data = 8'h04;
    16'h019A: data = 8'h80;
    16'h01A6: data = 8'h20;
    16'h01AD: data = 8'h01;
    16'h01AE: data = 8'h20;
    16'h01B1: data = 8'h02;
    16'h01B2: data = 8'h20;
    16'h01C1: data = 8'h05;
    16'h01C2: data = 8'h80;
    16'h01CA: data = 8'h40;
    16'h01CD: data = 8'h01;
    16'h01CE: data = 8'h40;
    16'h01D1: data = 8'h01;
    16'h01D2: data = 8'h80;
    16'h01D5: data = 8'h02;
    16'h01D6: data = 8'h40;
    16'h01D9: data = 8'h03;
    16'h01DA: data = 8'h20;
    16'h01E5: data = 8'h04;
    16'h01E6: data = 8'h40;
    16'h01EA: data = 8'h80;
    16'h01ED: data = 8'h04;
    16'h01EE: data = 8'h20;
    16'h01F1: data = 8'h14;
    16'h01F2: data = 8'h40;
    16'h01F5: data = 8'h02;
    16'h01F6: data = 8'h80;
    16'h0445: data = 8'h07;
    16'h0446: data = 8'h02;
    16'h0447: data = 8'h10;
    16'h0451: data = 8'h08;
    16'h0452: data = 8'h01;
    16'h0453: data = 8'h08;
    16'h049D: data = 8'h06;
    16'h049E: data = 8'h80;
    16'h0529: data = 8'h14;
    16'h052A: data = 8'h20;
    16'h0569: data = 8'h06;
    16'h056A: data = 8'h01;
    16'h05AD: data = 8'h08;
    16'h05AE: data = 8'h08;
    16'h05C9: data = 8'h08;
    16'h05CA: data = 8'h04;
    16'h05D1: data = 8'h08;
    16'h05D2: data = 8'h10;
    16'h05D5: data = 8'h08;
    16'h05D6: data = 8'h02;
    16'h0835: data = 8'h03;
    16'h0836: data = 8'h40;
    16'h0838: data = 8'h70;
    16'h0839: data = 8'h27;
    16'h083A: data = 8'h80;
    16'h0846: data = 8'h01;
    16'h0847: data = 8'h10;
    16'h084B: data = 8'h04;
    16'h0851: data = 8'h08;
    16'h0852: data = 8'h01;
    16'h0853: data = 8'h08;
    16'h0855: data = 8'h12;
    16'h0856: data = 8'h01;
    16'h0859: data = 8'h13;
    16'h085A: data = 8'h01;
    16'h0869: data = 8'h10;
    16'h086A: data = 8'h02;
    16'h086D: data = 8'h11;
    16'h086E: data = 8'h02;
    16'h0871: data = 8'h11;
    16'h0872: data = 8'h01;
    16'h0875: data = 8'h12;
    16'h0876: data = 8'h02;
    16'h0879: data = 8'h05;
    16'h087A: data = 8'h40;
    16'h0885: data = 8'h10;
    16'h0886: data = 8'h08;
    16'h0889: data = 8'h10;
    16'h088A: data = 8'h04;
    16'h088D: data = 8'h11;
    16'h088E: data = 8'h04;
    16'h0891: data = 8'h12;
    16'h0892: data = 8'h04;
    16'h0895: data = 8'h13;
    16'h0896: data = 8'h08;
    16'h0899: data = 8'h13;
    16'h089A: data = 8'h04;
    16'h08A5: data = 8'h07;
    16'h08A6: data = 8'h01;
    16'h08A9: data = 8'h10;
    16'h08AA: data = 8'h10;
    16'h08AD: data = 8'h11;
    16'h08AE: data = 8'h08;
    16'h08B1: data = 8'h12;
    16'h08B2: data = 8'h10;
    16'h08B5: data = 8'h12;
    16'h08B6: data = 8'h08;
    16'h08B9: data = 8'h13;
    16'h08BA: data = 8'h10;
    16'h08C5: data = 8'h17;
    16'h08C6: data = 8'h08;
    16'h08C9: data = 8'h17;
    16'h08CA: data = 8'h10;
    16'h08CD: data = 8'h16;
    16'h08CE: data = 8'h10;
    16'h08D1: data = 8'h11;
    16'h08D2: data = 8'h10;
    16'h08D5: data = 8'h15;
    16'h08D6: data = 8'h10;
    16'h08D9: data = 8'h14;
    16'h08DA: data = 8'h10;
    16'h08E9: data = 8'h17;
    16'h08EA: data = 8'h04;
    16'h08ED: data = 8'h16;
    16'h08EE: data = 8'h08;
    16'h08F1: data = 8'h15;
    16'h08F2: data = 8'h08;
    16'h08F5: data = 8'h14;
    16'h08F6: data = 8'h20;
    16'h08F9: data = 8'h14;
    16'h08FA: data = 8'h04;
    16'h0905: data = 8'h06;
    16'h0906: data = 8'h20;
    16'h0909: data = 8'h16;
    16'h090A: data = 8'h04;
    16'h090D: data = 8'h15;
    16'h090E: data = 8'h04;
    16'h0911: data = 8'h15;
    16'h0912: data = 8'h02;
    16'h0915: data = 8'h05;
    16'h0916: data = 8'h20;
    16'h0919: data = 8'h14;
    16'h091A: data = 8'h02;
    16'h0925: data = 8'h06;
    16'h0926: data = 8'h40;
    16'h0929: data = 8'h15;
    16'h092A: data = 8'h20;
    16'h092D: data = 8'h16;
    16'h092E: data = 8'h02;
    16'h0935: data = 8'h15;
    16'h0936: data = 8'h01;
    16'h0938: data = 8'h70;
    16'h0939: data = 8'h20;
    16'h093A: data = 8'h04;
    16'h0948: data = 8'h70;
    16'h0949: data = 8'h21;
    16'h094A: data = 8'h08;
    16'h0950: data = 8'h70;
    16'h0951: data = 8'h26;
    16'h0952: data = 8'h10;
    16'h0961: data = 8'h03;
    16'h0962: data = 8'h80;
    16'h0967: data = 8'h04;
    16'h0969: data = 8'h06;
    16'h096A: data = 8'h01;
    16'h096D: data = 8'h14;
    16'h096E: data = 8'h40;
    16'h0975: data = 8'h15;
    16'h0976: data = 8'h40;
    16'h0984: data = 8'h70;
    16'h0985: data = 8'h22;
    16'h0986: data = 8'h02;
    16'h09A6: data = 8'h20;
    16'h09AD: data = 8'h01;
    16'h09AE: data = 8'h20;
    16'h09B1: data = 8'h02;
    16'h09B2: data = 8'h20;
    16'h09C1: data = 8'h05;
    16'h09C2: data = 8'h80;
    16'h09CA: data = 8'h40;
    16'h09CD: data = 8'h01;
    16'h09CE: data = 8'h40;
    16'h09D1: data = 8'h01;
    16'h09D2: data = 8'h80;
    16'h09D5: data = 8'h02;
    16'h09D6: data = 8'h40;
    16'h09D9: data = 8'h03;
    16'h09DA: data = 8'h20;
    16'h09E5: data = 8'h04;
    16'h09E6: data = 8'h40;
    16'h09EA: data = 8'h80;
    16'h09ED: data = 8'h04;
    16'h09EE: data = 8'h20;
    16'h09F1: data = 8'h14;
    16'h09F2: data = 8'h40;
    16'h09F5: data = 8'h02;
    16'h09F6: data = 8'h80;
    16'h0C45: data = 8'h07;
    16'h0C46: data = 8'h02;
    16'h0C47: data = 8'h10;
    16'h0C51: data = 8'h08;
    16'h0C52: data = 8'h01;
    16'h0C53: data = 8'h08;
    16'h0C9D: data = 8'h06;
    16'h0C9E: data = 8'h80;
    16'h0D29: data = 8'h14;
    16'h0D2A: data = 8'h20;
    16'h0D69: data = 8'h06;
    16'h0D6A: data = 8'h01;
    16'h0DAD: data = 8'h08;
    16'h0DAE: data = 8'h08;
    16'h0DC9: data = 8'h08;
    16'h0DCA: data = 8'h04;
    16'h0DD1: data = 8'h08;
    16'h0DD2: data = 8'h10;
    16'h0DD5: data = 8'h08;
    16'h0DD6: data = 8'h02;
    16'h1035: data = 8'h03;
    16'h1036: data = 8'h40;
    16'h1046: data = 8'h01;
    16'h1047: data = 8'h10;
    16'h104B: data = 8'h04;
    16'h1051: data = 8'h08;
    16'h1052: data = 8'h01;
    16'h1053: data = 8'h08;
    16'h10A5: data = 8'h07;
    16'h10A6: data = 8'h01;
    16'h1161: data = 8'h03;
    16'h1162: data = 8'h80;
    16'h1167: data = 8'h04;
    16'h1169: data = 8'h06;
    16'h116A: data = 8'h01;
    16'h11A6: data = 8'h20;
    16'h11AD: data = 8'h01;
    16'h11AE: data = 8'h20;
    16'h11B1: data = 8'h02;
    16'h11B2: data = 8'h20;
    16'h11C1: data = 8'h05;
    16'h11C2: data = 8'h80;
    16'h11CA: data = 8'h40;
    16'h11CD: data = 8'h01;
    16'h11CE: data = 8'h40;
    16'h11D1: data = 8'h01;
    16'h11D2: data = 8'h80;
    16'h11D5: data = 8'h02;
    16'h11D6: data = 8'h40;
    16'h11D9: data = 8'h03;
    16'h11DA: data = 8'h20;
    16'h11E5: data = 8'h04;
    16'h11E6: data = 8'h40;
    16'h11EA: data = 8'h80;
    16'h11ED: data = 8'h04;
    16'h11EE: data = 8'h20;
    16'h11F1: data = 8'h14;
    16'h11F2: data = 8'h40;
    16'h11F5: data = 8'h02;
    16'h11F6: data = 8'h80;
    16'h1445: data = 8'h07;
    16'h1446: data = 8'h02;
    16'h1447: data = 8'h10;
    16'h1451: data = 8'h08;
    16'h1452: data = 8'h01;
    16'h1453: data = 8'h08;
    16'h149D: data = 8'h06;
    16'h149E: data = 8'h80;
    16'h1529: data = 8'h14;
    16'h152A: data = 8'h20;
    16'h1569: data = 8'h06;
    16'h156A: data = 8'h01;
    16'h15AD: data = 8'h08;
    16'h15AE: data = 8'h08;
    16'h15C9: data = 8'h08;
    16'h15CA: data = 8'h04;
    16'h15D1: data = 8'h08;
    16'h15D2: data = 8'h10;
    16'h15D5: data = 8'h08;
    16'h15D6: data = 8'h02;
    16'h1835: data = 8'h03;
    16'h1836: data = 8'h40;
    16'h1846: data = 8'h01;
    16'h1847: data = 8'h10;
    16'h184B: data = 8'h04;
    16'h1851: data = 8'h08;
    16'h1852: data = 8'h01;
    16'h1853: data = 8'h08;
    16'h18A5: data = 8'h07;
    16'h18A6: data = 8'h01;
    16'h1961: data = 8'h03;
    16'h1962: data = 8'h80;
    16'h1967: data = 8'h04;
    16'h1969: data = 8'h06;
    16'h196A: data = 8'h01;
    16'h19A6: data = 8'h20;
    16'h19AD: data = 8'h01;
    16'h19AE: data = 8'h20;
    16'h19B1: data = 8'h02;
    16'h19B2: data = 8'h20;
    16'h19C1: data = 8'h05;
    16'h19C2: data = 8'h80;
    16'h19CA: data = 8'h40;
    16'h19CD: data = 8'h01;
    16'h19CE: data = 8'h40;
    16'h19D1: data = 8'h01;
    16'h19D2: data = 8'h80;
    16'h19D5: data = 8'h02;
    16'h19D6: data = 8'h40;
    16'h19D9: data = 8'h03;
    16'h19DA: data = 8'h20;
    16'h19E5: data = 8'h04;
    16'h19E6: data = 8'h40;
    16'h19EA: data = 8'h80;
    16'h19ED: data = 8'h04;
    16'h19EE: data = 8'h20;
    16'h19F1: data = 8'h14;
    16'h19F2: data = 8'h40;
    16'h19F5: data = 8'h02;
    16'h19F6: data = 8'h80;
    16'h1C45: data = 8'h07;
    16'h1C46: data = 8'h02;
    16'h1C47: data = 8'h10;
    16'h1C51: data = 8'h08;
    16'h1C52: data = 8'h01;
    16'h1C53: data = 8'h08;
    16'h1C9D: data = 8'h06;
    16'h1C9E: data = 8'h80;
    16'h1D29: data = 8'h14;
    16'h1D2A: data = 8'h20;
    16'h1D69: data = 8'h06;
    16'h1D6A: data = 8'h01;
    16'h1DAD: data = 8'h08;
    16'h1DAE: data = 8'h08;
    16'h1DC9: data = 8'h08;
    16'h1DCA: data = 8'h04;
    16'h1DD1: data = 8'h08;
    16'h1DD2: data = 8'h10;
    16'h1DD5: data = 8'h08;
    16'h1DD6: data = 8'h02;
    16'h2035: data = 8'h03;
    16'h2036: data = 8'h40;
    16'h2046: data = 8'h01;
    16'h2047: data = 8'h10;
    16'h204B: data = 8'h04;
    16'h2051: data = 8'h08;
    16'h2052: data = 8'h01;
    16'h2053: data = 8'h08;
    16'h20A5: data = 8'h07;
    16'h20A6: data = 8'h01;
    16'h2161: data = 8'h03;
    16'h2162: data = 8'h80;
    16'h2167: data = 8'h04;
    16'h2169: data = 8'h06;
    16'h216A: data = 8'h01;
    16'h21A6: data = 8'h20;
    16'h21AD: data = 8'h01;
    16'h21AE: data = 8'h20;
    16'h21B1: data = 8'h02;
    16'h21B2: data = 8'h20;
    16'h21C1: data = 8'h05;
    16'h21C2: data = 8'h80;
    16'h21CA: data = 8'h40;
    16'h21CD: data = 8'h01;
    16'h21CE: data = 8'h40;
    16'h21D1: data = 8'h01;
    16'h21D2: data = 8'h80;
    16'h21D5: data = 8'h02;
    16'h21D6: data = 8'h40;
    16'h21D9: data = 8'h03;
    16'h21DA: data = 8'h20;
    16'h21E5: data = 8'h04;
    16'h21E6: data = 8'h40;
    16'h21EA: data = 8'h80;
    16'h21ED: data = 8'h04;
    16'h21EE: data = 8'h20;
    16'h21F1: data = 8'h14;
    16'h21F2: data = 8'h40;
    16'h21F5: data = 8'h02;
    16'h21F6: data = 8'h80;
    16'h2445: data = 8'h07;
    16'h2446: data = 8'h02;
    16'h2447: data = 8'h10;
    16'h2451: data = 8'h08;
    16'h2452: data = 8'h01;
    16'h2453: data = 8'h08;
    16'h249D: data = 8'h06;
    16'h249E: data = 8'h80;
    16'h2529: data = 8'h14;
    16'h252A: data = 8'h20;
    16'h2569: data = 8'h06;
    16'h256A: data = 8'h01;
    16'h25AD: data = 8'h08;
    16'h25AE: data = 8'h08;
    16'h25C9: data = 8'h08;
    16'h25CA: data = 8'h04;
    16'h25D1: data = 8'h08;
    16'h25D2: data = 8'h10;
    16'h25D5: data = 8'h08;
    16'h25D6: data = 8'h02;
    16'h2835: data = 8'h03;
    16'h2836: data = 8'h40;
    16'h2846: data = 8'h01;
    16'h2847: data = 8'h10;
    16'h284B: data = 8'h04;
    16'h2851: data = 8'h08;
    16'h2852: data = 8'h01;
    16'h2853: data = 8'h08;
    16'h28A5: data = 8'h07;
    16'h28A6: data = 8'h01;
    16'h2961: data = 8'h03;
    16'h2962: data = 8'h80;
    16'h2967: data = 8'h04;
    16'h2969: data = 8'h06;
    16'h296A: data = 8'h01;
    16'h29A6: data = 8'h20;
    16'h29AD: data = 8'h01;
    16'h29AE: data = 8'h20;
    16'h29B1: data = 8'h02;
    16'h29B2: data = 8'h20;
    16'h29C1: data = 8'h05;
    16'h29C2: data = 8'h80;
    16'h29CA: data = 8'h40;
    16'h29CD: data = 8'h01;
    16'h29CE: data = 8'h40;
    16'h29D1: data = 8'h01;
    16'h29D2: data = 8'h80;
    16'h29D5: data = 8'h02;
    16'h29D6: data = 8'h40;
    16'h29D9: data = 8'h03;
    16'h29DA: data = 8'h20;
    16'h29E5: data = 8'h04;
    16'h29E6: data = 8'h40;
    16'h29EA: data = 8'h80;
    16'h29ED: data = 8'h04;
    16'h29EE: data = 8'h20;
    16'h29F1: data = 8'h14;
    16'h29F2: data = 8'h40;
    16'h29F5: data = 8'h02;
    16'h29F6: data = 8'h80;
    16'h2C45: data = 8'h07;
    16'h2C46: data = 8'h02;
    16'h2C47: data = 8'h10;
    16'h2C51: data = 8'h08;
    16'h2C52: data = 8'h01;
    16'h2C53: data = 8'h08;
    16'h2C9D: data = 8'h06;
    16'h2C9E: data = 8'h80;
    16'h2D29: data = 8'h14;
    16'h2D2A: data = 8'h20;
    16'h2D69: data = 8'h06;
    16'h2D6A: data = 8'h01;
    16'h2DAD: data = 8'h08;
    16'h2DAE: data = 8'h08;
    16'h2DC9: data = 8'h08;
    16'h2DCA: data = 8'h04;
    16'h2DD1: data = 8'h08;
    16'h2DD2: data = 8'h10;
    16'h2DD5: data = 8'h08;
    16'h2DD6: data = 8'h02;
    16'h300F: data = 8'h20;
    16'h3035: data = 8'h03;
    16'h3036: data = 8'h40;
    16'h3046: data = 8'h01;
    16'h3047: data = 8'h10;
    16'h304B: data = 8'h04;
    16'h3051: data = 8'h08;
    16'h3052: data = 8'h01;
    16'h3053: data = 8'h08;
    16'h30A5: data = 8'h07;
    16'h30A6: data = 8'h01;
    16'h3161: data = 8'h03;
    16'h3162: data = 8'h80;
    16'h3167: data = 8'h04;
    16'h3169: data = 8'h06;
    16'h316A: data = 8'h01;
    16'h319B: data = 8'h80;
    16'h31A6: data = 8'h20;
    16'h31AD: data = 8'h01;
    16'h31AE: data = 8'h20;
    16'h31B1: data = 8'h02;
    16'h31B2: data = 8'h20;
    16'h31C1: data = 8'h05;
    16'h31C2: data = 8'h80;
    16'h31C7: data = 8'h40;
    16'h31CA: data = 8'h40;
    16'h31CD: data = 8'h01;
    16'h31CE: data = 8'h40;
    16'h31D1: data = 8'h01;
    16'h31D2: data = 8'h80;
    16'h31D5: data = 8'h02;
    16'h31D6: data = 8'h40;
    16'h31D9: data = 8'h03;
    16'h31DA: data = 8'h20;
    16'h31E5: data = 8'h04;
    16'h31E6: data = 8'h40;
    16'h31EA: data = 8'h80;
    16'h31ED: data = 8'h04;
    16'h31EE: data = 8'h20;
    16'h31F1: data = 8'h14;
    16'h31F2: data = 8'h40;
    16'h31F5: data = 8'h02;
    16'h31F6: data = 8'h80;
    16'h3445: data = 8'h07;
    16'h3446: data = 8'h02;
    16'h3447: data = 8'h10;
    16'h3451: data = 8'h08;
    16'h3452: data = 8'h01;
    16'h3453: data = 8'h08;
    16'h349D: data = 8'h06;
    16'h349E: data = 8'h80;
    16'h3529: data = 8'h14;
    16'h352A: data = 8'h20;
    16'h3569: data = 8'h06;
    16'h356A: data = 8'h01;
    16'h35AD: data = 8'h08;
    16'h35AE: data = 8'h08;
    16'h35C7: data = 8'h40;
    16'h35C9: data = 8'h08;
    16'h35CA: data = 8'h04;
    16'h35D1: data = 8'h08;
    16'h35D2: data = 8'h10;
    16'h35D5: data = 8'h08;
    16'h35D6: data = 8'h02;
    16'h3835: data = 8'h03;
    16'h3836: data = 8'h40;
    16'h3846: data = 8'h01;
    16'h3847: data = 8'h10;
    16'h384B: data = 8'h04;
    16'h3851: data = 8'h08;
    16'h3852: data = 8'h01;
    16'h3853: data = 8'h08;
    16'h38A5: data = 8'h07;
    16'h38A6: data = 8'h01;
    16'h3961: data = 8'h03;
    16'h3962: data = 8'h80;
    16'h3967: data = 8'h04;
    16'h3969: data = 8'h06;
    16'h396A: data = 8'h01;
    16'h39A6: data = 8'h20;
    16'h39AD: data = 8'h01;
    16'h39AE: data = 8'h20;
    16'h39B1: data = 8'h02;
    16'h39B2: data = 8'h20;
    16'h39C1: data = 8'h05;
    16'h39C2: data = 8'h80;
    16'h39CA: data = 8'h40;
    16'h39CD: data = 8'h01;
    16'h39CE: data = 8'h40;
    16'h39D1: data = 8'h01;
    16'h39D2: data = 8'h80;
    16'h39D5: data = 8'h02;
    16'h39D6: data = 8'h40;
    16'h39D9: data = 8'h03;
    16'h39DA: data = 8'h20;
    16'h39E5: data = 8'h04;
    16'h39E6: data = 8'h40;
    16'h39EA: data = 8'h80;
    16'h39ED: data = 8'h04;
    16'h39EE: data = 8'h20;
    16'h39F1: data = 8'h14;
    16'h39F2: data = 8'h40;
    16'h39F5: data = 8'h02;
    16'h39F6: data = 8'h80;
    16'h3C45: data = 8'h07;
    16'h3C46: data = 8'h02;
    16'h3C47: data = 8'h10;
    16'h3C51: data = 8'h08;
    16'h3C52: data = 8'h01;
    16'h3C53: data = 8'h08;
    16'h3C9D: data = 8'h06;
    16'h3C9E: data = 8'h80;
    16'h3D29: data = 8'h14;
    16'h3D2A: data = 8'h20;
    16'h3D69: data = 8'h06;
    16'h3D6A: data = 8'h01;
    16'h3DAD: data = 8'h08;
    16'h3DAE: data = 8'h08;
    16'h3DC9: data = 8'h08;
    16'h3DCA: data = 8'h04;
    16'h3DD1: data = 8'h08;
    16'h3DD2: data = 8'h10;
    16'h3DD5: data = 8'h08;
    16'h3DD6: data = 8'h02;
    default: data = 8'h00;
  endcase;
end

endmodule
