-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80ef",
     9 => x"b8080b0b",
    10 => x"80efbc08",
    11 => x"0b0b80ef",
    12 => x"c0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"efc00c0b",
    16 => x"0b80efbc",
    17 => x"0c0b0b80",
    18 => x"efb80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80e5c8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80efb870",
    57 => x"81f08827",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c5188ea",
    62 => x"04820b0b",
    63 => x"0b80ead8",
    64 => x"0c800b80",
    65 => x"efd00c80",
    66 => x"0b80efc8",
    67 => x"0c800b80",
    68 => x"efcc0c04",
    69 => x"02fc050d",
    70 => x"f880518f",
    71 => x"0b80efc8",
    72 => x"0c9f0b80",
    73 => x"efcc0ca0",
    74 => x"71708105",
    75 => x"533480ef",
    76 => x"cc08ff05",
    77 => x"80efcc0c",
    78 => x"80efcc08",
    79 => x"8025e838",
    80 => x"80efc808",
    81 => x"ff0580ef",
    82 => x"c80c80ef",
    83 => x"c8088025",
    84 => x"d038800b",
    85 => x"80efcc0c",
    86 => x"800b80ef",
    87 => x"c80c0284",
    88 => x"050d0402",
    89 => x"f0050df8",
    90 => x"8053f8a0",
    91 => x"5483bf52",
    92 => x"73708105",
    93 => x"55335170",
    94 => x"73708105",
    95 => x"5534ff12",
    96 => x"52718025",
    97 => x"eb38fbc0",
    98 => x"539f52a0",
    99 => x"73708105",
   100 => x"5534ff12",
   101 => x"52718025",
   102 => x"f2380290",
   103 => x"050d0402",
   104 => x"f4050d74",
   105 => x"538e0b80",
   106 => x"efc80825",
   107 => x"913882e3",
   108 => x"2d80efc8",
   109 => x"08ff0580",
   110 => x"efc80c83",
   111 => x"a50480ef",
   112 => x"c80880ef",
   113 => x"cc085351",
   114 => x"728a2e09",
   115 => x"8106be38",
   116 => x"7151719f",
   117 => x"24a43880",
   118 => x"efc808a0",
   119 => x"2911f880",
   120 => x"115151a0",
   121 => x"713480ef",
   122 => x"cc088105",
   123 => x"80efcc0c",
   124 => x"80efcc08",
   125 => x"519f7125",
   126 => x"de38800b",
   127 => x"80efcc0c",
   128 => x"80efc808",
   129 => x"810580ef",
   130 => x"c80c84a3",
   131 => x"0470a029",
   132 => x"12f88011",
   133 => x"51517271",
   134 => x"3480efcc",
   135 => x"08810580",
   136 => x"efcc0c80",
   137 => x"efcc08a0",
   138 => x"2e098106",
   139 => x"9138800b",
   140 => x"80efcc0c",
   141 => x"80efc808",
   142 => x"810580ef",
   143 => x"c80c028c",
   144 => x"050d0402",
   145 => x"e8050d77",
   146 => x"79565688",
   147 => x"0bfc1677",
   148 => x"712c8f06",
   149 => x"54525480",
   150 => x"53727225",
   151 => x"95387153",
   152 => x"fbe01451",
   153 => x"87713481",
   154 => x"14ff1454",
   155 => x"5472f138",
   156 => x"7153f915",
   157 => x"76712c87",
   158 => x"06535171",
   159 => x"802e8b38",
   160 => x"fbe01451",
   161 => x"71713481",
   162 => x"1454728e",
   163 => x"2495388f",
   164 => x"733153fb",
   165 => x"e01451a0",
   166 => x"71348114",
   167 => x"ff145454",
   168 => x"72f13802",
   169 => x"98050d04",
   170 => x"02f4050d",
   171 => x"800b80ef",
   172 => x"d00cf68c",
   173 => x"08f69008",
   174 => x"71882c72",
   175 => x"81ff0653",
   176 => x"54545171",
   177 => x"71258738",
   178 => x"820b80ef",
   179 => x"d00c7288",
   180 => x"2c7381ff",
   181 => x"06525271",
   182 => x"71258b38",
   183 => x"80efd008",
   184 => x"840780ef",
   185 => x"d00c820b",
   186 => x"0b0b80ea",
   187 => x"d80c830b",
   188 => x"f6880cfc",
   189 => x"0880efd0",
   190 => x"08515174",
   191 => x"802e8538",
   192 => x"70810751",
   193 => x"70f6940c",
   194 => x"feb80bf6",
   195 => x"800cff9c",
   196 => x"0bf6840c",
   197 => x"028c050d",
   198 => x"0402f405",
   199 => x"0d745372",
   200 => x"70810554",
   201 => x"80f52d52",
   202 => x"71802e89",
   203 => x"38715183",
   204 => x"9f2d869f",
   205 => x"04810b80",
   206 => x"efb80c02",
   207 => x"8c050d04",
   208 => x"02fc050d",
   209 => x"80e78c51",
   210 => x"86992d80",
   211 => x"e7bc51b7",
   212 => x"d02d80ef",
   213 => x"b808802e",
   214 => x"943880e7",
   215 => x"c45180c4",
   216 => x"842d80e7",
   217 => x"d05180c4",
   218 => x"842d86f4",
   219 => x"0480e7e0",
   220 => x"5186992d",
   221 => x"0284050d",
   222 => x"0402f005",
   223 => x"0d765375",
   224 => x"5280ec9c",
   225 => x"0b80f52d",
   226 => x"5180d2f9",
   227 => x"2d80efb8",
   228 => x"085480ef",
   229 => x"b808802e",
   230 => x"883880eb",
   231 => x"805187a5",
   232 => x"0480ebf8",
   233 => x"5190e52d",
   234 => x"7380efb8",
   235 => x"0c029005",
   236 => x"0d0402fc",
   237 => x"050d800b",
   238 => x"80ec9c0b",
   239 => x"81b72d86",
   240 => x"f95180c3",
   241 => x"db2d7251",
   242 => x"80c3b62d",
   243 => x"0284050d",
   244 => x"0402fc05",
   245 => x"0d810b80",
   246 => x"ec9c0b81",
   247 => x"b72d86f9",
   248 => x"5180c3db",
   249 => x"2d725180",
   250 => x"c3b62d02",
   251 => x"84050d04",
   252 => x"02cc050d",
   253 => x"800b80e7",
   254 => x"fc530298",
   255 => x"05705355",
   256 => x"5580c8b5",
   257 => x"2d735202",
   258 => x"a4055388",
   259 => x"9b047452",
   260 => x"81157452",
   261 => x"5580c988",
   262 => x"2d735272",
   263 => x"5180c8b5",
   264 => x"2d80e884",
   265 => x"52725180",
   266 => x"c8d72d72",
   267 => x"51b9962d",
   268 => x"80efb808",
   269 => x"d93880e8",
   270 => x"8c518699",
   271 => x"2d725186",
   272 => x"992d80e8",
   273 => x"fc518699",
   274 => x"2d725180",
   275 => x"e2d22d80",
   276 => x"efb80880",
   277 => x"2e883880",
   278 => x"eb805188",
   279 => x"e20480eb",
   280 => x"f85190e5",
   281 => x"2d02b405",
   282 => x"0d0402f0",
   283 => x"050df008",
   284 => x"8106538a",
   285 => x"fc2d8cf2",
   286 => x"2d8faa2d",
   287 => x"9ea62d81",
   288 => x"f92d7285",
   289 => x"38850bec",
   290 => x"0c8f8f2d",
   291 => x"8aa12d82",
   292 => x"942d8151",
   293 => x"85a82d84",
   294 => x"0bec0c80",
   295 => x"e89c5186",
   296 => x"992da18d",
   297 => x"2d80efb8",
   298 => x"08802e80",
   299 => x"db387284",
   300 => x"3886c02d",
   301 => x"80d5b52d",
   302 => x"80eadc51",
   303 => x"90e52d80",
   304 => x"5185a82d",
   305 => x"840bec0c",
   306 => x"8bb32d90",
   307 => x"f82d80ef",
   308 => x"b8085380",
   309 => x"d1d82d80",
   310 => x"ecf008fc",
   311 => x"0c80ecf0",
   312 => x"08862a81",
   313 => x"06528051",
   314 => x"80d2a32d",
   315 => x"80ecf008",
   316 => x"872a8106",
   317 => x"52815180",
   318 => x"d2a32d86",
   319 => x"54728338",
   320 => x"845473ec",
   321 => x"0c89c804",
   322 => x"800b80ef",
   323 => x"b80c0290",
   324 => x"050d0480",
   325 => x"0bffb00c",
   326 => x"04ffb008",
   327 => x"80efb80c",
   328 => x"04810bff",
   329 => x"b00c0402",
   330 => x"f8050d8a",
   331 => x"932d8a99",
   332 => x"2d80efb8",
   333 => x"0880efd4",
   334 => x"0880efb8",
   335 => x"083280ef",
   336 => x"d40c80ef",
   337 => x"b8088106",
   338 => x"52527080",
   339 => x"2e8d3880",
   340 => x"eca00851",
   341 => x"70802e83",
   342 => x"38702d71",
   343 => x"812a7081",
   344 => x"06515170",
   345 => x"802e8d38",
   346 => x"80eca408",
   347 => x"5170802e",
   348 => x"8338702d",
   349 => x"8aa12d02",
   350 => x"88050d04",
   351 => x"02fc050d",
   352 => x"80eca051",
   353 => x"80717084",
   354 => x"05530c80",
   355 => x"710c0284",
   356 => x"050d0402",
   357 => x"fc050d72",
   358 => x"8aa70b98",
   359 => x"0c517081",
   360 => x"248c3870",
   361 => x"842980ec",
   362 => x"a0057471",
   363 => x"0c510284",
   364 => x"050d0402",
   365 => x"f4050d80",
   366 => x"efd8518e",
   367 => x"992d80ef",
   368 => x"b8085280",
   369 => x"efb80880",
   370 => x"2e819d38",
   371 => x"8cd60480",
   372 => x"efb80881",
   373 => x"f02e0981",
   374 => x"068a3881",
   375 => x"0b80ece8",
   376 => x"0c8cd604",
   377 => x"80efb808",
   378 => x"81e02e09",
   379 => x"81068a38",
   380 => x"810b80ec",
   381 => x"ec0c8cd6",
   382 => x"0480efb8",
   383 => x"085280ec",
   384 => x"ec08802e",
   385 => x"893880ef",
   386 => x"b8088180",
   387 => x"05527184",
   388 => x"2c728f06",
   389 => x"535380ec",
   390 => x"e808802e",
   391 => x"9a387284",
   392 => x"2980eca8",
   393 => x"05721381",
   394 => x"712b7009",
   395 => x"73080673",
   396 => x"0c515353",
   397 => x"8cca0472",
   398 => x"842980ec",
   399 => x"a8057213",
   400 => x"83712b72",
   401 => x"0807720c",
   402 => x"5353800b",
   403 => x"80ecec0c",
   404 => x"800b80ec",
   405 => x"e80c80ef",
   406 => x"d8518dd4",
   407 => x"2d80efb8",
   408 => x"08ff24fe",
   409 => x"ea388052",
   410 => x"7180efb8",
   411 => x"0c028c05",
   412 => x"0d0402f8",
   413 => x"050d80ec",
   414 => x"a8528f51",
   415 => x"80727084",
   416 => x"05540cff",
   417 => x"11517080",
   418 => x"25f23802",
   419 => x"88050d04",
   420 => x"02f0050d",
   421 => x"7570822c",
   422 => x"fc0680ec",
   423 => x"a8117210",
   424 => x"9e067108",
   425 => x"70722a82",
   426 => x"732b7009",
   427 => x"7306750c",
   428 => x"53830680",
   429 => x"efb80c57",
   430 => x"53515351",
   431 => x"0290050d",
   432 => x"0402fc05",
   433 => x"0d725180",
   434 => x"710c800b",
   435 => x"84120c02",
   436 => x"84050d04",
   437 => x"02f0050d",
   438 => x"75700884",
   439 => x"12085353",
   440 => x"53ff5471",
   441 => x"712ea838",
   442 => x"8a932d84",
   443 => x"13087084",
   444 => x"29148811",
   445 => x"70087081",
   446 => x"ff068418",
   447 => x"08811187",
   448 => x"06841a0c",
   449 => x"53515551",
   450 => x"51518aa1",
   451 => x"2d715473",
   452 => x"80efb80c",
   453 => x"0290050d",
   454 => x"0402f405",
   455 => x"0d747008",
   456 => x"84120853",
   457 => x"53537072",
   458 => x"248f3872",
   459 => x"08841408",
   460 => x"71713152",
   461 => x"52528ec6",
   462 => x"04720884",
   463 => x"14087171",
   464 => x"31880552",
   465 => x"52527180",
   466 => x"efb80c02",
   467 => x"8c050d04",
   468 => x"02f8050d",
   469 => x"e008708b",
   470 => x"2a708106",
   471 => x"51525270",
   472 => x"802ea138",
   473 => x"80efd808",
   474 => x"70842980",
   475 => x"efe00573",
   476 => x"81ff0671",
   477 => x"0c515180",
   478 => x"efd80881",
   479 => x"11870680",
   480 => x"efd80c51",
   481 => x"800b80f0",
   482 => x"800c0288",
   483 => x"050d0402",
   484 => x"f8050d80",
   485 => x"efd8518d",
   486 => x"c12d8cf2",
   487 => x"2d8ed052",
   488 => x"80518b93",
   489 => x"2d028805",
   490 => x"0d04800b",
   491 => x"80ecf40c",
   492 => x"81c60b80",
   493 => x"ecf00c04",
   494 => x"80f08408",
   495 => x"80efb80c",
   496 => x"0402fc05",
   497 => x"0d8fcb04",
   498 => x"8bb32d87",
   499 => x"518d902d",
   500 => x"80efb808",
   501 => x"f33880da",
   502 => x"518d902d",
   503 => x"80efb808",
   504 => x"e73880ef",
   505 => x"b80880ec",
   506 => x"f40c80ef",
   507 => x"b8085185",
   508 => x"a82d0284",
   509 => x"050d0402",
   510 => x"f4050d80",
   511 => x"f0840853",
   512 => x"82942d80",
   513 => x"0b80f088",
   514 => x"0c720880",
   515 => x"2e80d138",
   516 => x"820b80ef",
   517 => x"cc0c80f0",
   518 => x"88088f06",
   519 => x"80efc80c",
   520 => x"7208812e",
   521 => x"098106a1",
   522 => x"3880ecf0",
   523 => x"08881408",
   524 => x"2c708106",
   525 => x"51527180",
   526 => x"2e883880",
   527 => x"e8b45190",
   528 => x"c60480e8",
   529 => x"b8518699",
   530 => x"2d841308",
   531 => x"5186992d",
   532 => x"80f08808",
   533 => x"810580f0",
   534 => x"880c8c13",
   535 => x"53908904",
   536 => x"028c050d",
   537 => x"047180f0",
   538 => x"840c8ff7",
   539 => x"2d80f088",
   540 => x"08ff0580",
   541 => x"f08c0c04",
   542 => x"02e8050d",
   543 => x"80f08408",
   544 => x"80f09008",
   545 => x"56568751",
   546 => x"8d902d80",
   547 => x"efb80881",
   548 => x"2a708106",
   549 => x"51527180",
   550 => x"2eac3891",
   551 => x"a1048bb3",
   552 => x"2d87518d",
   553 => x"902d80ef",
   554 => x"b808f338",
   555 => x"80ecf408",
   556 => x"81327080",
   557 => x"ecf40c51",
   558 => x"85a82d80",
   559 => x"ecf40880",
   560 => x"2e84388c",
   561 => x"f22d80ec",
   562 => x"f4087054",
   563 => x"5271802e",
   564 => x"84ce3881",
   565 => x"f5518d90",
   566 => x"2d80efb8",
   567 => x"08812a70",
   568 => x"81065152",
   569 => x"71802eb3",
   570 => x"3880f08c",
   571 => x"08527180",
   572 => x"2e8a38ff",
   573 => x"1280f08c",
   574 => x"0c929b04",
   575 => x"80f08808",
   576 => x"1080f088",
   577 => x"08057084",
   578 => x"29175152",
   579 => x"88120880",
   580 => x"2e8938ff",
   581 => x"51881208",
   582 => x"52712d81",
   583 => x"f2518d90",
   584 => x"2d80efb8",
   585 => x"08812a70",
   586 => x"81065152",
   587 => x"71802eb4",
   588 => x"3880f088",
   589 => x"08ff1180",
   590 => x"f08c0856",
   591 => x"53537372",
   592 => x"258a3881",
   593 => x"1480f08c",
   594 => x"0c92e404",
   595 => x"72101370",
   596 => x"84291751",
   597 => x"52881208",
   598 => x"802e8938",
   599 => x"fe518812",
   600 => x"0852712d",
   601 => x"81fd518d",
   602 => x"902d80ef",
   603 => x"b808812a",
   604 => x"70810651",
   605 => x"52719738",
   606 => x"81eb518d",
   607 => x"902d80ef",
   608 => x"b808812a",
   609 => x"70810651",
   610 => x"5271802e",
   611 => x"b13880f0",
   612 => x"8c08802e",
   613 => x"8a38800b",
   614 => x"80f08c0c",
   615 => x"93be0480",
   616 => x"f0880810",
   617 => x"80f08808",
   618 => x"05708429",
   619 => x"17515288",
   620 => x"1208802e",
   621 => x"8938fd51",
   622 => x"88120852",
   623 => x"712d81fa",
   624 => x"518d902d",
   625 => x"80efb808",
   626 => x"812a7081",
   627 => x"06515271",
   628 => x"973881f4",
   629 => x"518d902d",
   630 => x"80efb808",
   631 => x"812a7081",
   632 => x"06515271",
   633 => x"802eb138",
   634 => x"80f08808",
   635 => x"ff115452",
   636 => x"80f08c08",
   637 => x"73258938",
   638 => x"7280f08c",
   639 => x"0c949804",
   640 => x"71101270",
   641 => x"84291751",
   642 => x"52881208",
   643 => x"802e8938",
   644 => x"fc518812",
   645 => x"0852712d",
   646 => x"80f08c08",
   647 => x"70535473",
   648 => x"802e8738",
   649 => x"ff145494",
   650 => x"9f04820b",
   651 => x"80efcc0c",
   652 => x"718f0680",
   653 => x"efc80c80",
   654 => x"da518d90",
   655 => x"2d80efb8",
   656 => x"08812a70",
   657 => x"81065152",
   658 => x"71802e81",
   659 => x"8a3880f0",
   660 => x"840880f0",
   661 => x"8c085553",
   662 => x"73802e8a",
   663 => x"388c13ff",
   664 => x"15555394",
   665 => x"d8047208",
   666 => x"5271822e",
   667 => x"a1387182",
   668 => x"26893871",
   669 => x"812ea538",
   670 => x"95d70471",
   671 => x"842e0981",
   672 => x"0680d438",
   673 => x"88130851",
   674 => x"90e52d95",
   675 => x"d70480f0",
   676 => x"8c085188",
   677 => x"13085271",
   678 => x"2d95d704",
   679 => x"810b8814",
   680 => x"082b80ec",
   681 => x"f0083280",
   682 => x"ecf00c8f",
   683 => x"f72d95d7",
   684 => x"04740880",
   685 => x"2ea43874",
   686 => x"08518d90",
   687 => x"2d80efb8",
   688 => x"08810652",
   689 => x"71802e8c",
   690 => x"3880f08c",
   691 => x"08518415",
   692 => x"0852712d",
   693 => x"88155574",
   694 => x"d8388054",
   695 => x"800b80ef",
   696 => x"cc0c738f",
   697 => x"0680efc8",
   698 => x"0ca05273",
   699 => x"80f08c08",
   700 => x"2e098106",
   701 => x"993880f0",
   702 => x"8808ff05",
   703 => x"74327009",
   704 => x"81057072",
   705 => x"079f2a91",
   706 => x"71315151",
   707 => x"53537151",
   708 => x"839f2d81",
   709 => x"14548e74",
   710 => x"25c23880",
   711 => x"ecf40853",
   712 => x"7280efb8",
   713 => x"0c029805",
   714 => x"0d0402f4",
   715 => x"050dd452",
   716 => x"81ff720c",
   717 => x"71085381",
   718 => x"ff720c72",
   719 => x"882b83fe",
   720 => x"80067208",
   721 => x"7081ff06",
   722 => x"51525381",
   723 => x"ff720c72",
   724 => x"7107882b",
   725 => x"72087081",
   726 => x"ff065152",
   727 => x"5381ff72",
   728 => x"0c727107",
   729 => x"882b7208",
   730 => x"7081ff06",
   731 => x"720780ef",
   732 => x"b80c5253",
   733 => x"028c050d",
   734 => x"0402f405",
   735 => x"0d747671",
   736 => x"81ff06d4",
   737 => x"0c535380",
   738 => x"f0940885",
   739 => x"3871892b",
   740 => x"5271982a",
   741 => x"d40c7190",
   742 => x"2a7081ff",
   743 => x"06d40c51",
   744 => x"71882a70",
   745 => x"81ff06d4",
   746 => x"0c517181",
   747 => x"ff06d40c",
   748 => x"72902a70",
   749 => x"81ff06d4",
   750 => x"0c51d408",
   751 => x"7081ff06",
   752 => x"515182b8",
   753 => x"bf527081",
   754 => x"ff2e0981",
   755 => x"06943881",
   756 => x"ff0bd40c",
   757 => x"d4087081",
   758 => x"ff06ff14",
   759 => x"54515171",
   760 => x"e5387080",
   761 => x"efb80c02",
   762 => x"8c050d04",
   763 => x"02fc050d",
   764 => x"81c75181",
   765 => x"ff0bd40c",
   766 => x"ff115170",
   767 => x"8025f438",
   768 => x"0284050d",
   769 => x"0402f405",
   770 => x"0d81ff0b",
   771 => x"d40c9353",
   772 => x"805287fc",
   773 => x"80c15196",
   774 => x"f92d80ef",
   775 => x"b8088b38",
   776 => x"81ff0bd4",
   777 => x"0c815398",
   778 => x"b30497ec",
   779 => x"2dff1353",
   780 => x"72de3872",
   781 => x"80efb80c",
   782 => x"028c050d",
   783 => x"0402ec05",
   784 => x"0d810b80",
   785 => x"f0940c84",
   786 => x"54d00870",
   787 => x"8f2a7081",
   788 => x"06515153",
   789 => x"72f33872",
   790 => x"d00c97ec",
   791 => x"2d80e8bc",
   792 => x"5186992d",
   793 => x"d008708f",
   794 => x"2a708106",
   795 => x"51515372",
   796 => x"f338810b",
   797 => x"d00cb153",
   798 => x"805284d4",
   799 => x"80c05196",
   800 => x"f92d80ef",
   801 => x"b808812e",
   802 => x"93387282",
   803 => x"2ebf38ff",
   804 => x"135372e4",
   805 => x"38ff1454",
   806 => x"73ffae38",
   807 => x"97ec2d83",
   808 => x"aa52849c",
   809 => x"80c85196",
   810 => x"f92d80ef",
   811 => x"b808812e",
   812 => x"09810693",
   813 => x"3896aa2d",
   814 => x"80efb808",
   815 => x"83ffff06",
   816 => x"537283aa",
   817 => x"2e9f3898",
   818 => x"852d99e0",
   819 => x"0480e8c8",
   820 => x"5186992d",
   821 => x"80539bb5",
   822 => x"0480e8e0",
   823 => x"5186992d",
   824 => x"80549b86",
   825 => x"0481ff0b",
   826 => x"d40cb154",
   827 => x"97ec2d8f",
   828 => x"cf538052",
   829 => x"87fc80f7",
   830 => x"5196f92d",
   831 => x"80efb808",
   832 => x"5580efb8",
   833 => x"08812e09",
   834 => x"81069c38",
   835 => x"81ff0bd4",
   836 => x"0c820a52",
   837 => x"849c80e9",
   838 => x"5196f92d",
   839 => x"80efb808",
   840 => x"802e8d38",
   841 => x"97ec2dff",
   842 => x"135372c6",
   843 => x"389af904",
   844 => x"81ff0bd4",
   845 => x"0c80efb8",
   846 => x"085287fc",
   847 => x"80fa5196",
   848 => x"f92d80ef",
   849 => x"b808b238",
   850 => x"81ff0bd4",
   851 => x"0cd40853",
   852 => x"81ff0bd4",
   853 => x"0c81ff0b",
   854 => x"d40c81ff",
   855 => x"0bd40c81",
   856 => x"ff0bd40c",
   857 => x"72862a70",
   858 => x"81067656",
   859 => x"51537296",
   860 => x"3880efb8",
   861 => x"08549b86",
   862 => x"0473822e",
   863 => x"fedb38ff",
   864 => x"145473fe",
   865 => x"e7387380",
   866 => x"f0940c73",
   867 => x"8b388152",
   868 => x"87fc80d0",
   869 => x"5196f92d",
   870 => x"81ff0bd4",
   871 => x"0cd00870",
   872 => x"8f2a7081",
   873 => x"06515153",
   874 => x"72f33872",
   875 => x"d00c81ff",
   876 => x"0bd40c81",
   877 => x"537280ef",
   878 => x"b80c0294",
   879 => x"050d0402",
   880 => x"e8050d78",
   881 => x"5681ff0b",
   882 => x"d40cd008",
   883 => x"708f2a70",
   884 => x"81065151",
   885 => x"5372f338",
   886 => x"82810bd0",
   887 => x"0c81ff0b",
   888 => x"d40c7752",
   889 => x"87fc80d8",
   890 => x"5196f92d",
   891 => x"80efb808",
   892 => x"802e8d38",
   893 => x"80e8f051",
   894 => x"86992d81",
   895 => x"539cf804",
   896 => x"81ff0bd4",
   897 => x"0c81fe0b",
   898 => x"d40c80ff",
   899 => x"55757084",
   900 => x"05570870",
   901 => x"982ad40c",
   902 => x"70902c70",
   903 => x"81ff06d4",
   904 => x"0c547088",
   905 => x"2c7081ff",
   906 => x"06d40c54",
   907 => x"7081ff06",
   908 => x"d40c54ff",
   909 => x"15557480",
   910 => x"25d33881",
   911 => x"ff0bd40c",
   912 => x"81ff0bd4",
   913 => x"0c81ff0b",
   914 => x"d40c868d",
   915 => x"a05481ff",
   916 => x"0bd40cd4",
   917 => x"0881ff06",
   918 => x"55748738",
   919 => x"ff145473",
   920 => x"ed3881ff",
   921 => x"0bd40cd0",
   922 => x"08708f2a",
   923 => x"70810651",
   924 => x"515372f3",
   925 => x"3872d00c",
   926 => x"7280efb8",
   927 => x"0c029805",
   928 => x"0d0402e8",
   929 => x"050d7855",
   930 => x"805681ff",
   931 => x"0bd40cd0",
   932 => x"08708f2a",
   933 => x"70810651",
   934 => x"515372f3",
   935 => x"3882810b",
   936 => x"d00c81ff",
   937 => x"0bd40c77",
   938 => x"5287fc80",
   939 => x"d15196f9",
   940 => x"2d80dbc6",
   941 => x"df5480ef",
   942 => x"b808802e",
   943 => x"8b3880e9",
   944 => x"80518699",
   945 => x"2d9e9c04",
   946 => x"81ff0bd4",
   947 => x"0cd40870",
   948 => x"81ff0651",
   949 => x"537281fe",
   950 => x"2e098106",
   951 => x"9e3880ff",
   952 => x"5396aa2d",
   953 => x"80efb808",
   954 => x"75708405",
   955 => x"570cff13",
   956 => x"53728025",
   957 => x"ec388156",
   958 => x"9e8104ff",
   959 => x"145473c8",
   960 => x"3881ff0b",
   961 => x"d40c81ff",
   962 => x"0bd40cd0",
   963 => x"08708f2a",
   964 => x"70810651",
   965 => x"515372f3",
   966 => x"3872d00c",
   967 => x"7580efb8",
   968 => x"0c029805",
   969 => x"0d04800b",
   970 => x"80f6ac0c",
   971 => x"800b80f6",
   972 => x"b00c800b",
   973 => x"80f6a40c",
   974 => x"800b80f6",
   975 => x"b40c800b",
   976 => x"80f6b80c",
   977 => x"800b80f6",
   978 => x"bc0c800b",
   979 => x"80f6c00c",
   980 => x"800b80f6",
   981 => x"c40c800b",
   982 => x"80f6c80c",
   983 => x"800b80f6",
   984 => x"9c0c800b",
   985 => x"80f6a00c",
   986 => x"800b80f6",
   987 => x"cc0c800b",
   988 => x"80f6d00c",
   989 => x"800b80f6",
   990 => x"d40b818a",
   991 => x"2d820b80",
   992 => x"ed800c80",
   993 => x"0b80f6d8",
   994 => x"0c800b80",
   995 => x"f6dc0c80",
   996 => x"0b80f6e0",
   997 => x"0c800b80",
   998 => x"f6e40c80",
   999 => x"0b80f6a8",
  1000 => x"0c800b80",
  1001 => x"ecf80c04",
  1002 => x"02f8050d",
  1003 => x"735280f6",
  1004 => x"a408802e",
  1005 => x"94387182",
  1006 => x"2b83fc06",
  1007 => x"80f6e811",
  1008 => x"085252bd",
  1009 => x"ce2d9fda",
  1010 => x"04711083",
  1011 => x"fe0680f6",
  1012 => x"e81180e0",
  1013 => x"2d5252bd",
  1014 => x"f92d0288",
  1015 => x"050d0402",
  1016 => x"ec050d76",
  1017 => x"5574802e",
  1018 => x"80c5389a",
  1019 => x"1580e02d",
  1020 => x"51bdf92d",
  1021 => x"80efb808",
  1022 => x"80efb808",
  1023 => x"80f6dc0c",
  1024 => x"80efb808",
  1025 => x"545480f6",
  1026 => x"a408802e",
  1027 => x"9a389415",
  1028 => x"80e02d51",
  1029 => x"bdf92d80",
  1030 => x"efb80890",
  1031 => x"2b83fff0",
  1032 => x"0a067075",
  1033 => x"07515372",
  1034 => x"80f6dc0c",
  1035 => x"a0b40474",
  1036 => x"80f6dc0c",
  1037 => x"80f6dc08",
  1038 => x"5372802e",
  1039 => x"9d3880f6",
  1040 => x"9c08fe14",
  1041 => x"712980f6",
  1042 => x"b8080580",
  1043 => x"f6e00c70",
  1044 => x"842b80f6",
  1045 => x"a80c54a1",
  1046 => x"880480f6",
  1047 => x"bc0880f6",
  1048 => x"dc0c80f6",
  1049 => x"c00880f6",
  1050 => x"e00c80f6",
  1051 => x"a408802e",
  1052 => x"8b3880f6",
  1053 => x"9c08842b",
  1054 => x"53a18304",
  1055 => x"80f6c408",
  1056 => x"842b5372",
  1057 => x"80f6a80c",
  1058 => x"0294050d",
  1059 => x"0402d805",
  1060 => x"0d800b80",
  1061 => x"f6a40c84",
  1062 => x"5498bd2d",
  1063 => x"80efb808",
  1064 => x"802e9738",
  1065 => x"80f09852",
  1066 => x"80519d82",
  1067 => x"2d80efb8",
  1068 => x"08802e86",
  1069 => x"38fe54a1",
  1070 => x"c204ff14",
  1071 => x"54738024",
  1072 => x"d838738d",
  1073 => x"3880e990",
  1074 => x"5186992d",
  1075 => x"7355a8e1",
  1076 => x"04800b80",
  1077 => x"f6d80c81",
  1078 => x"0b80f6e4",
  1079 => x"0c885380",
  1080 => x"e9a45280",
  1081 => x"f0ce5180",
  1082 => x"ca862d80",
  1083 => x"efb80889",
  1084 => x"3880efb8",
  1085 => x"0880f6e4",
  1086 => x"0c885380",
  1087 => x"e9b05280",
  1088 => x"f0ea5180",
  1089 => x"ca862d80",
  1090 => x"efb80889",
  1091 => x"3880efb8",
  1092 => x"0880f6e4",
  1093 => x"0c80f6e4",
  1094 => x"08802e81",
  1095 => x"8c3880f3",
  1096 => x"de0b80f5",
  1097 => x"2d80f3df",
  1098 => x"0b80f52d",
  1099 => x"71982b71",
  1100 => x"902b0780",
  1101 => x"f3e00b80",
  1102 => x"f52d7088",
  1103 => x"2b720780",
  1104 => x"f3e10b80",
  1105 => x"f52d7107",
  1106 => x"7080f6d8",
  1107 => x"0c80f496",
  1108 => x"0b80f52d",
  1109 => x"80f4970b",
  1110 => x"80f52d71",
  1111 => x"882b0757",
  1112 => x"5f51525a",
  1113 => x"56575574",
  1114 => x"81abaa2e",
  1115 => x"09810691",
  1116 => x"387351bd",
  1117 => x"ce2d80ef",
  1118 => x"b80880f6",
  1119 => x"d80ca38f",
  1120 => x"047482d4",
  1121 => x"d52e8838",
  1122 => x"80e9bc51",
  1123 => x"a3e00480",
  1124 => x"f0985280",
  1125 => x"f6d80851",
  1126 => x"9d822d80",
  1127 => x"efb80855",
  1128 => x"80efb808",
  1129 => x"802e85b9",
  1130 => x"38885380",
  1131 => x"e9b05280",
  1132 => x"f0ea5180",
  1133 => x"ca862d80",
  1134 => x"efb8088a",
  1135 => x"38810b80",
  1136 => x"f6a40ca3",
  1137 => x"e6048853",
  1138 => x"80e9a452",
  1139 => x"80f0ce51",
  1140 => x"80ca862d",
  1141 => x"80efb808",
  1142 => x"802e8b38",
  1143 => x"80e9d051",
  1144 => x"86992da4",
  1145 => x"c50480f4",
  1146 => x"960b80f5",
  1147 => x"2d547380",
  1148 => x"d52e0981",
  1149 => x"0680ce38",
  1150 => x"80f4970b",
  1151 => x"80f52d54",
  1152 => x"7381aa2e",
  1153 => x"098106bd",
  1154 => x"38800b80",
  1155 => x"f0980b80",
  1156 => x"f52d5654",
  1157 => x"7481e92e",
  1158 => x"83388154",
  1159 => x"7481eb2e",
  1160 => x"8c388055",
  1161 => x"73752e09",
  1162 => x"810684b5",
  1163 => x"3880f0a3",
  1164 => x"0b80f52d",
  1165 => x"56758e38",
  1166 => x"80f0a40b",
  1167 => x"80f52d54",
  1168 => x"73822e86",
  1169 => x"388055a8",
  1170 => x"e10480f0",
  1171 => x"a50b80f5",
  1172 => x"2d7080f6",
  1173 => x"9c0cff05",
  1174 => x"7080f6a0",
  1175 => x"0c558176",
  1176 => x"80f6cc0c",
  1177 => x"70760655",
  1178 => x"5773802e",
  1179 => x"97387476",
  1180 => x"56588115",
  1181 => x"7710707a",
  1182 => x"06565855",
  1183 => x"73f43874",
  1184 => x"80f6cc0c",
  1185 => x"80f0a60b",
  1186 => x"80f52d80",
  1187 => x"f0a70b80",
  1188 => x"f52d5680",
  1189 => x"f6d80805",
  1190 => x"75828029",
  1191 => x"057080f6",
  1192 => x"b40c80f0",
  1193 => x"a80b80f5",
  1194 => x"2d7080f6",
  1195 => x"c80c80f6",
  1196 => x"a4085957",
  1197 => x"5876802e",
  1198 => x"82c83888",
  1199 => x"5380e9b0",
  1200 => x"5280f0ea",
  1201 => x"5180ca86",
  1202 => x"2d805580",
  1203 => x"efb80875",
  1204 => x"2e098106",
  1205 => x"838b3880",
  1206 => x"f69c0870",
  1207 => x"842b80f6",
  1208 => x"a80c7080",
  1209 => x"f6c40c80",
  1210 => x"f0bd0b80",
  1211 => x"f52d80f0",
  1212 => x"bc0b80f5",
  1213 => x"2d718280",
  1214 => x"290580f0",
  1215 => x"be0b80f5",
  1216 => x"2d708480",
  1217 => x"80291280",
  1218 => x"f0bf0b80",
  1219 => x"f52d7081",
  1220 => x"800a2912",
  1221 => x"7080f6d0",
  1222 => x"0c80f6c8",
  1223 => x"08712980",
  1224 => x"f6b40805",
  1225 => x"7080f6b8",
  1226 => x"0c80f0c5",
  1227 => x"0b80f52d",
  1228 => x"80f0c40b",
  1229 => x"80f52d71",
  1230 => x"82802905",
  1231 => x"80f0c60b",
  1232 => x"80f52d70",
  1233 => x"84808029",
  1234 => x"1280f0c7",
  1235 => x"0b80f52d",
  1236 => x"70982b81",
  1237 => x"f00a0672",
  1238 => x"057080f6",
  1239 => x"bc0c80f0",
  1240 => x"c90b80f5",
  1241 => x"2d80f0c8",
  1242 => x"0b80f52d",
  1243 => x"71882b07",
  1244 => x"57465257",
  1245 => x"52575d57",
  1246 => x"51525f52",
  1247 => x"5c575757",
  1248 => x"7580f6d4",
  1249 => x"0b818a2d",
  1250 => x"fe147729",
  1251 => x"750580f6",
  1252 => x"c00c820b",
  1253 => x"80ed800c",
  1254 => x"80f6a408",
  1255 => x"802e81ba",
  1256 => x"3880f098",
  1257 => x"5280f6d8",
  1258 => x"0816519d",
  1259 => x"822d80ef",
  1260 => x"b808802e",
  1261 => x"81a43884",
  1262 => x"5380e5d8",
  1263 => x"5280f494",
  1264 => x"5180ca86",
  1265 => x"2d80efb8",
  1266 => x"08818f38",
  1267 => x"80f4810b",
  1268 => x"80f52d80",
  1269 => x"f4800b80",
  1270 => x"f52d7188",
  1271 => x"2b0780f4",
  1272 => x"820b80f5",
  1273 => x"2d70902b",
  1274 => x"720780f4",
  1275 => x"830b80f5",
  1276 => x"2d70982b",
  1277 => x"720780ed",
  1278 => x"800c5b52",
  1279 => x"58555aa8",
  1280 => x"da0480f0",
  1281 => x"aa0b80f5",
  1282 => x"2d80f0a9",
  1283 => x"0b80f52d",
  1284 => x"71828029",
  1285 => x"057080f6",
  1286 => x"a80c70a0",
  1287 => x"2983ff05",
  1288 => x"70892a70",
  1289 => x"80f6c40c",
  1290 => x"80f0af0b",
  1291 => x"80f52d80",
  1292 => x"f0ae0b80",
  1293 => x"f52d7182",
  1294 => x"80290570",
  1295 => x"80f6d00c",
  1296 => x"7b71291e",
  1297 => x"7080f6c0",
  1298 => x"0c7d80f6",
  1299 => x"bc0c7305",
  1300 => x"80f6b80c",
  1301 => x"5a545151",
  1302 => x"55598051",
  1303 => x"9fdf2d81",
  1304 => x"557480ef",
  1305 => x"b80c02a8",
  1306 => x"050d0402",
  1307 => x"f0050d80",
  1308 => x"ecfc0853",
  1309 => x"72802580",
  1310 => x"c73872fe",
  1311 => x"0a065372",
  1312 => x"fe0a2eb1",
  1313 => x"38805480",
  1314 => x"f6c80874",
  1315 => x"2ea73880",
  1316 => x"f6e85280",
  1317 => x"ecfc08fe",
  1318 => x"0a0680f6",
  1319 => x"b4080574",
  1320 => x"80f6d008",
  1321 => x"2905519b",
  1322 => x"bf2d8114",
  1323 => x"5480f6c8",
  1324 => x"087426db",
  1325 => x"3880ecfc",
  1326 => x"08fe0a06",
  1327 => x"80ecfc0c",
  1328 => x"0290050d",
  1329 => x"0402f005",
  1330 => x"0d757087",
  1331 => x"2a555380",
  1332 => x"f6a40885",
  1333 => x"3872882a",
  1334 => x"5480ecfc",
  1335 => x"08fe0a06",
  1336 => x"5373732e",
  1337 => x"a338a8eb",
  1338 => x"2d80f6e8",
  1339 => x"5280f6b4",
  1340 => x"0814519d",
  1341 => x"822d80ef",
  1342 => x"b8085380",
  1343 => x"efb80880",
  1344 => x"2e883873",
  1345 => x"80ecfc0c",
  1346 => x"81537280",
  1347 => x"efb80c02",
  1348 => x"90050d04",
  1349 => x"02f4050d",
  1350 => x"74705253",
  1351 => x"a9c52d80",
  1352 => x"efb80852",
  1353 => x"80efb808",
  1354 => x"802e8b38",
  1355 => x"72519fa8",
  1356 => x"2d80efb8",
  1357 => x"08527180",
  1358 => x"efb80c02",
  1359 => x"8c050d04",
  1360 => x"02f8050d",
  1361 => x"73527151",
  1362 => x"a9c52d80",
  1363 => x"efb80889",
  1364 => x"3880efb8",
  1365 => x"0852aaec",
  1366 => x"0471519f",
  1367 => x"a82d80ef",
  1368 => x"b808802e",
  1369 => x"87388112",
  1370 => x"52aac604",
  1371 => x"7180efb8",
  1372 => x"0c028805",
  1373 => x"0d0402f4",
  1374 => x"050d7480",
  1375 => x"f6a40852",
  1376 => x"5370802e",
  1377 => x"9e388073",
  1378 => x"80ffffff",
  1379 => x"f8065252",
  1380 => x"7080ffff",
  1381 => x"fff82e09",
  1382 => x"81068338",
  1383 => x"81527151",
  1384 => x"abaf0472",
  1385 => x"83ffff2e",
  1386 => x"09810683",
  1387 => x"38815170",
  1388 => x"80efb80c",
  1389 => x"028c050d",
  1390 => x"0402f405",
  1391 => x"0d747671",
  1392 => x"535452a9",
  1393 => x"c52d80ef",
  1394 => x"b808802e",
  1395 => x"80c63880",
  1396 => x"f6a40880",
  1397 => x"2e9b3871",
  1398 => x"822b83fc",
  1399 => x"0680f6e8",
  1400 => x"11745351",
  1401 => x"52bdce2d",
  1402 => x"80efb808",
  1403 => x"720cac89",
  1404 => x"04711083",
  1405 => x"fe0680f6",
  1406 => x"e8117453",
  1407 => x"5152bdf9",
  1408 => x"2d80efb8",
  1409 => x"0872818a",
  1410 => x"2d80ecfc",
  1411 => x"08810a07",
  1412 => x"80ecfc0c",
  1413 => x"028c050d",
  1414 => x"0402dc05",
  1415 => x"0d7b80f6",
  1416 => x"9c088480",
  1417 => x"291cff11",
  1418 => x"892a7080",
  1419 => x"f6cc082a",
  1420 => x"705a5a51",
  1421 => x"5559fe0a",
  1422 => x"0b80ecfc",
  1423 => x"0c80ed80",
  1424 => x"0851aac0",
  1425 => x"2d80efb8",
  1426 => x"0880efb8",
  1427 => x"08595581",
  1428 => x"7725a038",
  1429 => x"811551aa",
  1430 => x"c02d80ef",
  1431 => x"b80880ef",
  1432 => x"b8085375",
  1433 => x"5254abb9",
  1434 => x"2d73ff17",
  1435 => x"57557581",
  1436 => x"24e238f0",
  1437 => x"0a5480f6",
  1438 => x"a4088538",
  1439 => x"83ffff54",
  1440 => x"73527451",
  1441 => x"abb92d78",
  1442 => x"802e8838",
  1443 => x"77527851",
  1444 => x"abb92da8",
  1445 => x"eb2d7609",
  1446 => x"81055580",
  1447 => x"f6a40880",
  1448 => x"2e81ab38",
  1449 => x"80f09852",
  1450 => x"80f6d40b",
  1451 => x"80e02d80",
  1452 => x"f6d80805",
  1453 => x"519d822d",
  1454 => x"80efb808",
  1455 => x"802e818e",
  1456 => x"38845380",
  1457 => x"e5d85280",
  1458 => x"f4945180",
  1459 => x"ca862d80",
  1460 => x"efb80880",
  1461 => x"f93880f4",
  1462 => x"810b80f5",
  1463 => x"2d80f480",
  1464 => x"0b80f52d",
  1465 => x"71882b07",
  1466 => x"80f4820b",
  1467 => x"80f52d70",
  1468 => x"902b7207",
  1469 => x"80f4830b",
  1470 => x"80f52d70",
  1471 => x"982b7207",
  1472 => x"7a115152",
  1473 => x"5b525255",
  1474 => x"567380f4",
  1475 => x"800b81b7",
  1476 => x"2d73882a",
  1477 => x"557480f4",
  1478 => x"810b81b7",
  1479 => x"2d73902a",
  1480 => x"557480f4",
  1481 => x"820b81b7",
  1482 => x"2d73982a",
  1483 => x"557480f4",
  1484 => x"830b81b7",
  1485 => x"2d7380ed",
  1486 => x"800c80f0",
  1487 => x"985280f6",
  1488 => x"d40b80e0",
  1489 => x"2d80f6d8",
  1490 => x"0805519b",
  1491 => x"bf2d7780",
  1492 => x"efb80c02",
  1493 => x"a4050d04",
  1494 => x"02ec050d",
  1495 => x"76558070",
  1496 => x"7680f52d",
  1497 => x"53545270",
  1498 => x"722e8338",
  1499 => x"81537081",
  1500 => x"e52e9f38",
  1501 => x"81707406",
  1502 => x"52547080",
  1503 => x"2e94388b",
  1504 => x"1580f52d",
  1505 => x"70832a70",
  1506 => x"76065152",
  1507 => x"55708338",
  1508 => x"73527180",
  1509 => x"efb80c02",
  1510 => x"94050d04",
  1511 => x"02e4050d",
  1512 => x"7970842c",
  1513 => x"1a718f06",
  1514 => x"52555372",
  1515 => x"8a3880f0",
  1516 => x"98527351",
  1517 => x"9d822d72",
  1518 => x"a02980f0",
  1519 => x"98055480",
  1520 => x"7480f52d",
  1521 => x"56537473",
  1522 => x"2e833881",
  1523 => x"537481e5",
  1524 => x"2e81f138",
  1525 => x"72802e81",
  1526 => x"eb388b14",
  1527 => x"80f52d70",
  1528 => x"832a8106",
  1529 => x"58567699",
  1530 => x"3880ecf8",
  1531 => x"08537289",
  1532 => x"387280f4",
  1533 => x"980b81b7",
  1534 => x"2d7680ec",
  1535 => x"f80cb1c4",
  1536 => x"04758f2e",
  1537 => x"09810681",
  1538 => x"bb38749f",
  1539 => x"068d2980",
  1540 => x"f48b1151",
  1541 => x"53811480",
  1542 => x"f52d7370",
  1543 => x"81055581",
  1544 => x"b72d8314",
  1545 => x"80f52d73",
  1546 => x"70810555",
  1547 => x"81b72d85",
  1548 => x"1480f52d",
  1549 => x"73708105",
  1550 => x"5581b72d",
  1551 => x"871480f5",
  1552 => x"2d737081",
  1553 => x"055581b7",
  1554 => x"2d891480",
  1555 => x"f52d7370",
  1556 => x"81055581",
  1557 => x"b72d8e14",
  1558 => x"80f52d73",
  1559 => x"70810555",
  1560 => x"81b72d90",
  1561 => x"1480f52d",
  1562 => x"73708105",
  1563 => x"5581b72d",
  1564 => x"921480f5",
  1565 => x"2d737081",
  1566 => x"055581b7",
  1567 => x"2d941480",
  1568 => x"f52d7370",
  1569 => x"81055581",
  1570 => x"b72d9614",
  1571 => x"80f52d73",
  1572 => x"70810555",
  1573 => x"81b72d98",
  1574 => x"1480f52d",
  1575 => x"73708105",
  1576 => x"5581b72d",
  1577 => x"9c1480f5",
  1578 => x"2d737081",
  1579 => x"055581b7",
  1580 => x"2d9e1480",
  1581 => x"f52d7381",
  1582 => x"b72d80ec",
  1583 => x"f8088105",
  1584 => x"80ecf80c",
  1585 => x"7380efb8",
  1586 => x"0c029c05",
  1587 => x"0d0402e0",
  1588 => x"050d797b",
  1589 => x"59578070",
  1590 => x"5752b29b",
  1591 => x"0473ae2e",
  1592 => x"09810694",
  1593 => x"38718724",
  1594 => x"af387612",
  1595 => x"51a07181",
  1596 => x"b72d8112",
  1597 => x"52b1e504",
  1598 => x"76125572",
  1599 => x"8113ff9f",
  1600 => x"157081ff",
  1601 => x"06515353",
  1602 => x"54709926",
  1603 => x"86387281",
  1604 => x"df065473",
  1605 => x"7581b72d",
  1606 => x"81165680",
  1607 => x"76197080",
  1608 => x"f52d7081",
  1609 => x"ff065755",
  1610 => x"52557375",
  1611 => x"2e833881",
  1612 => x"55718a24",
  1613 => x"983874ff",
  1614 => x"a438718a",
  1615 => x"248f3876",
  1616 => x"1251a071",
  1617 => x"81b72d81",
  1618 => x"1252b2ba",
  1619 => x"04800b8b",
  1620 => x"1881b72d",
  1621 => x"02a0050d",
  1622 => x"0402ec05",
  1623 => x"0d76789c",
  1624 => x"11085355",
  1625 => x"55bdce2d",
  1626 => x"80efb808",
  1627 => x"84160c9a",
  1628 => x"1480e02d",
  1629 => x"51bdf92d",
  1630 => x"80efb808",
  1631 => x"80efb808",
  1632 => x"88170c80",
  1633 => x"efb80853",
  1634 => x"5380f6a4",
  1635 => x"08802e99",
  1636 => x"38941480",
  1637 => x"e02d51bd",
  1638 => x"f92d80ef",
  1639 => x"b808902b",
  1640 => x"83fff00a",
  1641 => x"06701451",
  1642 => x"52718816",
  1643 => x"0c80750c",
  1644 => x"810b80ef",
  1645 => x"b80c0294",
  1646 => x"050d0402",
  1647 => x"f4050d74",
  1648 => x"70088105",
  1649 => x"710c7008",
  1650 => x"80f6a008",
  1651 => x"06535371",
  1652 => x"8f388813",
  1653 => x"0851aa94",
  1654 => x"2d80efb8",
  1655 => x"0888140c",
  1656 => x"810b80ef",
  1657 => x"b80c028c",
  1658 => x"050d0402",
  1659 => x"f0050d75",
  1660 => x"881108fe",
  1661 => x"0580f69c",
  1662 => x"082980f6",
  1663 => x"b8080571",
  1664 => x"0880f6a0",
  1665 => x"08060580",
  1666 => x"efb80c54",
  1667 => x"0290050d",
  1668 => x"0402f805",
  1669 => x"0d7351b3",
  1670 => x"eb2d7452",
  1671 => x"80efb808",
  1672 => x"519d822d",
  1673 => x"0288050d",
  1674 => x"0402f005",
  1675 => x"0d758811",
  1676 => x"08fe0580",
  1677 => x"f69c0829",
  1678 => x"80f6b808",
  1679 => x"11720880",
  1680 => x"f6a00806",
  1681 => x"05795553",
  1682 => x"54549bbf",
  1683 => x"2d029005",
  1684 => x"0d0402ff",
  1685 => x"bc050d62",
  1686 => x"6466686a",
  1687 => x"4343435a",
  1688 => x"5a807071",
  1689 => x"72415e5e",
  1690 => x"5b7980f6",
  1691 => x"bc082e09",
  1692 => x"81068938",
  1693 => x"80f6a408",
  1694 => x"7b2e8338",
  1695 => x"815e8057",
  1696 => x"80f6a808",
  1697 => x"772e8193",
  1698 => x"38765278",
  1699 => x"51af9c2d",
  1700 => x"80efb808",
  1701 => x"567e9138",
  1702 => x"80efb808",
  1703 => x"51aed82d",
  1704 => x"80efb808",
  1705 => x"802ebb38",
  1706 => x"7c55761b",
  1707 => x"5480f498",
  1708 => x"53755260",
  1709 => x"517f2d80",
  1710 => x"efb80880",
  1711 => x"25863881",
  1712 => x"5cb5e204",
  1713 => x"800b80ef",
  1714 => x"b8082596",
  1715 => x"387b802e",
  1716 => x"80c93880",
  1717 => x"f0985276",
  1718 => x"842c1951",
  1719 => x"9bbf2db6",
  1720 => x"9b0480ec",
  1721 => x"f8085d80",
  1722 => x"778f0657",
  1723 => x"58758f2e",
  1724 => x"09810683",
  1725 => x"3881587b",
  1726 => x"802e9438",
  1727 => x"77802e8f",
  1728 => x"3880f098",
  1729 => x"5276842c",
  1730 => x"19519bbf",
  1731 => x"2d805c81",
  1732 => x"175780f6",
  1733 => x"a8087726",
  1734 => x"feef3880",
  1735 => x"f6a80877",
  1736 => x"26b4387d",
  1737 => x"802eaf38",
  1738 => x"7951aa94",
  1739 => x"2d80efb8",
  1740 => x"0880efb8",
  1741 => x"08525aaa",
  1742 => x"f62d80ef",
  1743 => x"b8089738",
  1744 => x"fe1a80f6",
  1745 => x"9c082980",
  1746 => x"f6b80805",
  1747 => x"80f6a808",
  1748 => x"1c5c59b4",
  1749 => x"fe040280",
  1750 => x"c4050d04",
  1751 => x"02ec050d",
  1752 => x"78557754",
  1753 => x"765380f6",
  1754 => x"e0085280",
  1755 => x"f6dc0851",
  1756 => x"b4d22d02",
  1757 => x"94050d04",
  1758 => x"02e8050d",
  1759 => x"77797c58",
  1760 => x"56547480",
  1761 => x"2ebe3888",
  1762 => x"53841452",
  1763 => x"745180ca",
  1764 => x"862d80ef",
  1765 => x"b808ad38",
  1766 => x"83538c14",
  1767 => x"52881551",
  1768 => x"80ca862d",
  1769 => x"80efb808",
  1770 => x"9b388174",
  1771 => x"0c749415",
  1772 => x"0c757c31",
  1773 => x"98150c75",
  1774 => x"9c150c79",
  1775 => x"90150c81",
  1776 => x"54b7c604",
  1777 => x"80547380",
  1778 => x"efb80c02",
  1779 => x"98050d04",
  1780 => x"02d0050d",
  1781 => x"80557d52",
  1782 => x"02b005e4",
  1783 => x"0551b1ce",
  1784 => x"2d8053b6",
  1785 => x"f85202b0",
  1786 => x"05e00551",
  1787 => x"b6dc2d74",
  1788 => x"802e8638",
  1789 => x"79519fdf",
  1790 => x"2d7480ef",
  1791 => x"b80c02b0",
  1792 => x"050d0402",
  1793 => x"cc050d80",
  1794 => x"567f5202",
  1795 => x"b405e405",
  1796 => x"51b1ce2d",
  1797 => x"8053b6f8",
  1798 => x"5202b405",
  1799 => x"e00551b6",
  1800 => x"dc2d7570",
  1801 => x"56547380",
  1802 => x"2e8d387a",
  1803 => x"527e51b2",
  1804 => x"d92d80ef",
  1805 => x"b8085574",
  1806 => x"80efb80c",
  1807 => x"02b4050d",
  1808 => x"0402c805",
  1809 => x"0d606053",
  1810 => x"02bc05e4",
  1811 => x"055256b1",
  1812 => x"ce2d8057",
  1813 => x"8053b6f8",
  1814 => x"5202b805",
  1815 => x"e00551b6",
  1816 => x"dc2d7580",
  1817 => x"2ea6387b",
  1818 => x"941180e0",
  1819 => x"2d5254bd",
  1820 => x"f92d80ef",
  1821 => x"b808902b",
  1822 => x"7c9a1180",
  1823 => x"e02d5355",
  1824 => x"55bdf92d",
  1825 => x"7480efb8",
  1826 => x"0807760c",
  1827 => x"7680efb8",
  1828 => x"0c02b805",
  1829 => x"0d0402f8",
  1830 => x"050d8052",
  1831 => x"7351b8c1",
  1832 => x"2d028805",
  1833 => x"0d0402f8",
  1834 => x"050d8075",
  1835 => x"7080f52d",
  1836 => x"51525270",
  1837 => x"81e52e09",
  1838 => x"81068338",
  1839 => x"81527009",
  1840 => x"81057080",
  1841 => x"25730770",
  1842 => x"54515170",
  1843 => x"802e8838",
  1844 => x"7377710c",
  1845 => x"51815271",
  1846 => x"80efb80c",
  1847 => x"0288050d",
  1848 => x"0402e005",
  1849 => x"0d797b9c",
  1850 => x"12085758",
  1851 => x"58815674",
  1852 => x"81aa3874",
  1853 => x"7780f52d",
  1854 => x"55567381",
  1855 => x"e52e0981",
  1856 => x"06833881",
  1857 => x"56730981",
  1858 => x"05708025",
  1859 => x"77077058",
  1860 => x"51547380",
  1861 => x"2e818538",
  1862 => x"88538418",
  1863 => x"52765180",
  1864 => x"c7de2d83",
  1865 => x"538c1852",
  1866 => x"88175180",
  1867 => x"c7de2d98",
  1868 => x"1880f52d",
  1869 => x"8b1881b7",
  1870 => x"2d748c18",
  1871 => x"81b72d74",
  1872 => x"8d1881b7",
  1873 => x"2d749618",
  1874 => x"818a2d74",
  1875 => x"8e18818a",
  1876 => x"2d749818",
  1877 => x"818a2d74",
  1878 => x"9018818a",
  1879 => x"2d749218",
  1880 => x"818a2d96",
  1881 => x"1880e02d",
  1882 => x"51bdf92d",
  1883 => x"80efb808",
  1884 => x"9a18818a",
  1885 => x"2d941880",
  1886 => x"e02d51bd",
  1887 => x"f92d80ef",
  1888 => x"b8089418",
  1889 => x"818a2d90",
  1890 => x"180851bd",
  1891 => x"ce2d80ef",
  1892 => x"b8089c18",
  1893 => x"0c810b9c",
  1894 => x"190cff56",
  1895 => x"7580efb8",
  1896 => x"0c02a005",
  1897 => x"0d0402c0",
  1898 => x"050d6163",
  1899 => x"71535957",
  1900 => x"b9962d80",
  1901 => x"5480efb8",
  1902 => x"08742e09",
  1903 => x"810681e6",
  1904 => x"38bbcc04",
  1905 => x"80efb808",
  1906 => x"54bc9d04",
  1907 => x"ff598153",
  1908 => x"b9a65202",
  1909 => x"a0057052",
  1910 => x"56b6dc2d",
  1911 => x"78802581",
  1912 => x"8a3880f6",
  1913 => x"a408802e",
  1914 => x"81813880",
  1915 => x"f6dc0854",
  1916 => x"7351a9c5",
  1917 => x"2d80efb8",
  1918 => x"08802ec8",
  1919 => x"3873519f",
  1920 => x"a82d80ef",
  1921 => x"b80851aa",
  1922 => x"f62d80ef",
  1923 => x"b8088e38",
  1924 => x"73519fa8",
  1925 => x"2d80efb8",
  1926 => x"0854bbf0",
  1927 => x"04735281",
  1928 => x"51ac992d",
  1929 => x"80efb808",
  1930 => x"fe0580f6",
  1931 => x"9c082980",
  1932 => x"f6b80805",
  1933 => x"55848053",
  1934 => x"805280f0",
  1935 => x"985180c8",
  1936 => x"892d8054",
  1937 => x"80f69c08",
  1938 => x"742e9638",
  1939 => x"80f09852",
  1940 => x"7315519b",
  1941 => x"bf2d8114",
  1942 => x"5480f69c",
  1943 => x"087426ec",
  1944 => x"388153b9",
  1945 => x"a6527551",
  1946 => x"b6dc2d80",
  1947 => x"54737924",
  1948 => x"b5387652",
  1949 => x"0280c005",
  1950 => x"e40551b1",
  1951 => x"ce2d775d",
  1952 => x"80527751",
  1953 => x"ac992d80",
  1954 => x"efb8085e",
  1955 => x"8040a002",
  1956 => x"bc0581b7",
  1957 => x"2d8153b9",
  1958 => x"e1520280",
  1959 => x"c005e005",
  1960 => x"51b6dc2d",
  1961 => x"7f547380",
  1962 => x"efb80c02",
  1963 => x"80c0050d",
  1964 => x"0402f405",
  1965 => x"0d80f6d0",
  1966 => x"0880f69c",
  1967 => x"0829872b",
  1968 => x"80f6c008",
  1969 => x"0580efb8",
  1970 => x"0c028c05",
  1971 => x"0d0402f4",
  1972 => x"050d7470",
  1973 => x"882a83fe",
  1974 => x"80067072",
  1975 => x"982a0772",
  1976 => x"882b87fc",
  1977 => x"80800671",
  1978 => x"0773982b",
  1979 => x"0780efb8",
  1980 => x"0c515351",
  1981 => x"028c050d",
  1982 => x"0402f805",
  1983 => x"0d028e05",
  1984 => x"80f52d74",
  1985 => x"882b0770",
  1986 => x"83ffff06",
  1987 => x"80efb80c",
  1988 => x"51028805",
  1989 => x"0d0402f4",
  1990 => x"050d7476",
  1991 => x"78535452",
  1992 => x"80712597",
  1993 => x"38727081",
  1994 => x"055480f5",
  1995 => x"2d727081",
  1996 => x"055481b7",
  1997 => x"2dff1151",
  1998 => x"70eb3880",
  1999 => x"7281b72d",
  2000 => x"028c050d",
  2001 => x"0402dc05",
  2002 => x"0d7a7c71",
  2003 => x"08565a56",
  2004 => x"73802e89",
  2005 => x"38ff1476",
  2006 => x"0c80c0b0",
  2007 => x"04841608",
  2008 => x"55815474",
  2009 => x"8b2481ca",
  2010 => x"388b1980",
  2011 => x"f52d7084",
  2012 => x"2a708106",
  2013 => x"771080f4",
  2014 => x"980b80f5",
  2015 => x"2d5c5351",
  2016 => x"55577380",
  2017 => x"2e80e738",
  2018 => x"7417822b",
  2019 => x"80c2de0b",
  2020 => x"80ed8c12",
  2021 => x"0c548416",
  2022 => x"08902984",
  2023 => x"17083170",
  2024 => x"1080faec",
  2025 => x"05515490",
  2026 => x"7481b72d",
  2027 => x"84160890",
  2028 => x"29841708",
  2029 => x"31701080",
  2030 => x"faed0551",
  2031 => x"54a07481",
  2032 => x"b72d7781",
  2033 => x"ff068417",
  2034 => x"08565473",
  2035 => x"802e8a38",
  2036 => x"9c5380f4",
  2037 => x"9852bfdd",
  2038 => x"048b5378",
  2039 => x"52749029",
  2040 => x"75317010",
  2041 => x"80faee05",
  2042 => x"525480c0",
  2043 => x"a5047417",
  2044 => x"822b80c0",
  2045 => x"dd0b80ed",
  2046 => x"8c120c54",
  2047 => x"7781ff06",
  2048 => x"84170856",
  2049 => x"5473802e",
  2050 => x"8b389c53",
  2051 => x"80f49852",
  2052 => x"80c09804",
  2053 => x"8b537852",
  2054 => x"74902975",
  2055 => x"31701080",
  2056 => x"faec0552",
  2057 => x"54841608",
  2058 => x"81058417",
  2059 => x"0cbe962d",
  2060 => x"80547380",
  2061 => x"efb80c02",
  2062 => x"a4050d04",
  2063 => x"02e8050d",
  2064 => x"77558056",
  2065 => x"805380c3",
  2066 => x"8e520298",
  2067 => x"05f80551",
  2068 => x"b6dc2d75",
  2069 => x"80efb80c",
  2070 => x"0298050d",
  2071 => x"0402ec05",
  2072 => x"0d80eeb8",
  2073 => x"08175180",
  2074 => x"c0bc2d80",
  2075 => x"efb80855",
  2076 => x"80efb808",
  2077 => x"802ea138",
  2078 => x"8b5380ef",
  2079 => x"b8085280",
  2080 => x"f49851be",
  2081 => x"962d80fa",
  2082 => x"e8085473",
  2083 => x"802e8938",
  2084 => x"745280f4",
  2085 => x"9851732d",
  2086 => x"0294050d",
  2087 => x"0402e005",
  2088 => x"0d80eeb8",
  2089 => x"08578058",
  2090 => x"8053bec5",
  2091 => x"5202a005",
  2092 => x"f80551b6",
  2093 => x"dc2d7755",
  2094 => x"748b24a2",
  2095 => x"38749029",
  2096 => x"75317010",
  2097 => x"80faec05",
  2098 => x"57548076",
  2099 => x"81b72d9e",
  2100 => x"16811670",
  2101 => x"5755568b",
  2102 => x"7425ef38",
  2103 => x"735802a0",
  2104 => x"050d0402",
  2105 => x"fc050d72",
  2106 => x"5170fd2e",
  2107 => x"b23870fd",
  2108 => x"248b3870",
  2109 => x"fc2e80d0",
  2110 => x"3880c2d2",
  2111 => x"0470fe2e",
  2112 => x"b93870ff",
  2113 => x"2e098106",
  2114 => x"80c83880",
  2115 => x"eeb80851",
  2116 => x"70802ebe",
  2117 => x"38ff1180",
  2118 => x"eeb80c80",
  2119 => x"c2d20480",
  2120 => x"eeb808f4",
  2121 => x"057080ee",
  2122 => x"b80c5170",
  2123 => x"8025a338",
  2124 => x"800b80ee",
  2125 => x"b80c80c2",
  2126 => x"d20480ee",
  2127 => x"b8088105",
  2128 => x"80eeb80c",
  2129 => x"80c2d204",
  2130 => x"80eeb808",
  2131 => x"8c0580ee",
  2132 => x"b80c80c1",
  2133 => x"9d2d8ff7",
  2134 => x"2d028405",
  2135 => x"0d0402fc",
  2136 => x"050d80ee",
  2137 => x"b8081351",
  2138 => x"80c0bc2d",
  2139 => x"80efb808",
  2140 => x"802e8938",
  2141 => x"80efb808",
  2142 => x"519fdf2d",
  2143 => x"800b80ee",
  2144 => x"b80c80c1",
  2145 => x"9d2d8ff7",
  2146 => x"2d028405",
  2147 => x"0d0402f4",
  2148 => x"050d7452",
  2149 => x"80720852",
  2150 => x"5370732e",
  2151 => x"8938ff11",
  2152 => x"720c80c3",
  2153 => x"ac047584",
  2154 => x"130c8153",
  2155 => x"7280efb8",
  2156 => x"0c028c05",
  2157 => x"0d0402fc",
  2158 => x"050d800b",
  2159 => x"80eeb80c",
  2160 => x"80c19d2d",
  2161 => x"8fb82d80",
  2162 => x"efb80880",
  2163 => x"eea80c80",
  2164 => x"ed845190",
  2165 => x"e52d0284",
  2166 => x"050d0471",
  2167 => x"80fae80c",
  2168 => x"0402f805",
  2169 => x"0dff1451",
  2170 => x"80527072",
  2171 => x"2e8b3881",
  2172 => x"1271812c",
  2173 => x"525270f7",
  2174 => x"38f71280",
  2175 => x"efb80c02",
  2176 => x"88050d04",
  2177 => x"02cc050d",
  2178 => x"8057840b",
  2179 => x"ec0c76fb",
  2180 => x"0c7e5202",
  2181 => x"a4057052",
  2182 => x"53b1ce2d",
  2183 => x"725280fd",
  2184 => x"f451b883",
  2185 => x"2d80efb8",
  2186 => x"08772e80",
  2187 => x"ec3880fd",
  2188 => x"f8087771",
  2189 => x"53595580",
  2190 => x"c3e12d80",
  2191 => x"efb80859",
  2192 => x"81577775",
  2193 => x"2580d238",
  2194 => x"78527751",
  2195 => x"84c32d80",
  2196 => x"f0985280",
  2197 => x"fdf451b4",
  2198 => x"912d80ef",
  2199 => x"b808802e",
  2200 => x"9c3880f0",
  2201 => x"985683fc",
  2202 => x"54757084",
  2203 => x"055708e8",
  2204 => x"0cfc1454",
  2205 => x"738025f1",
  2206 => x"3880c585",
  2207 => x"0480efb8",
  2208 => x"08578480",
  2209 => x"5580fdf4",
  2210 => x"51b3bb2d",
  2211 => x"fc801581",
  2212 => x"19595574",
  2213 => x"8024ffb0",
  2214 => x"3880fdf8",
  2215 => x"08f80c76",
  2216 => x"80efb80c",
  2217 => x"02b4050d",
  2218 => x"0402c405",
  2219 => x"0d606264",
  2220 => x"72545659",
  2221 => x"55b9962d",
  2222 => x"805380ef",
  2223 => x"b808732e",
  2224 => x"09810681",
  2225 => x"8c387352",
  2226 => x"7451bba6",
  2227 => x"2d80efb8",
  2228 => x"085380ef",
  2229 => x"b808802e",
  2230 => x"80f73881",
  2231 => x"5377802e",
  2232 => x"80ef3880",
  2233 => x"74525680",
  2234 => x"c3e12d80",
  2235 => x"efb80875",
  2236 => x"5302a405",
  2237 => x"70535457",
  2238 => x"b1ce2d72",
  2239 => x"5202bc05",
  2240 => x"f40551b8",
  2241 => x"832d80ef",
  2242 => x"b8085380",
  2243 => x"efb80876",
  2244 => x"2ebf3875",
  2245 => x"7425b838",
  2246 => x"76527551",
  2247 => x"84c32d80",
  2248 => x"f0985177",
  2249 => x"2d80efb8",
  2250 => x"08802e8e",
  2251 => x"3880f098",
  2252 => x"5202bc05",
  2253 => x"f40551b4",
  2254 => x"a92d02bc",
  2255 => x"05f40551",
  2256 => x"b3bb2dfc",
  2257 => x"80148117",
  2258 => x"57547380",
  2259 => x"24ca3881",
  2260 => x"537280ef",
  2261 => x"b80c02bc",
  2262 => x"050d0402",
  2263 => x"c8050d60",
  2264 => x"6202b405",
  2265 => x"56585372",
  2266 => x"802e8c38",
  2267 => x"72527351",
  2268 => x"b2d92d80",
  2269 => x"c789047f",
  2270 => x"52029c05",
  2271 => x"705253b1",
  2272 => x"ce2d7252",
  2273 => x"7351b883",
  2274 => x"2d80efb8",
  2275 => x"085480ef",
  2276 => x"b808802e",
  2277 => x"bf387c54",
  2278 => x"80745255",
  2279 => x"80c3e12d",
  2280 => x"80efb808",
  2281 => x"56747425",
  2282 => x"a9387552",
  2283 => x"745184c3",
  2284 => x"2d02ac05",
  2285 => x"705253b3",
  2286 => x"eb2d80ef",
  2287 => x"b8085176",
  2288 => x"2d7251b3",
  2289 => x"bb2dfc80",
  2290 => x"14811656",
  2291 => x"54738024",
  2292 => x"d9387c54",
  2293 => x"7380efb8",
  2294 => x"0c02b805",
  2295 => x"0d0402e8",
  2296 => x"050d7779",
  2297 => x"7b565656",
  2298 => x"80537274",
  2299 => x"25963872",
  2300 => x"16731652",
  2301 => x"527080f5",
  2302 => x"2d7281b7",
  2303 => x"2d811353",
  2304 => x"80c7ea04",
  2305 => x"0298050d",
  2306 => x"0402ec05",
  2307 => x"0d767902",
  2308 => x"88059f05",
  2309 => x"80f52d55",
  2310 => x"55558052",
  2311 => x"71742590",
  2312 => x"38711551",
  2313 => x"727181b7",
  2314 => x"2d811252",
  2315 => x"80c89c04",
  2316 => x"0294050d",
  2317 => x"0402f405",
  2318 => x"0d747653",
  2319 => x"53717081",
  2320 => x"055380f5",
  2321 => x"2d517073",
  2322 => x"70810555",
  2323 => x"81b72d70",
  2324 => x"ec38028c",
  2325 => x"050d0402",
  2326 => x"f4050d74",
  2327 => x"76545271",
  2328 => x"70810553",
  2329 => x"80f52d51",
  2330 => x"70f538ff",
  2331 => x"12527270",
  2332 => x"81055480",
  2333 => x"f52d5170",
  2334 => x"72708105",
  2335 => x"5481b72d",
  2336 => x"70ec3802",
  2337 => x"8c050d04",
  2338 => x"02d0050d",
  2339 => x"7d7f5859",
  2340 => x"885380df",
  2341 => x"5202a405",
  2342 => x"70525880",
  2343 => x"c8892d80",
  2344 => x"02b00581",
  2345 => x"b72d8756",
  2346 => x"7518778f",
  2347 => x"06555580",
  2348 => x"e9dc1480",
  2349 => x"f52d7581",
  2350 => x"b72d7684",
  2351 => x"2cff1757",
  2352 => x"57758424",
  2353 => x"e3388079",
  2354 => x"80f52d55",
  2355 => x"5673762e",
  2356 => x"a2387518",
  2357 => x"761a5555",
  2358 => x"7380f52d",
  2359 => x"7581b72d",
  2360 => x"81165675",
  2361 => x"84248c38",
  2362 => x"75197080",
  2363 => x"f52d5154",
  2364 => x"73e03889",
  2365 => x"5302b005",
  2366 => x"f4055278",
  2367 => x"5180c7de",
  2368 => x"2d02b005",
  2369 => x"0d0402e8",
  2370 => x"050d7779",
  2371 => x"7b585555",
  2372 => x"80537276",
  2373 => x"25a53874",
  2374 => x"70810556",
  2375 => x"80f52d74",
  2376 => x"70810556",
  2377 => x"80f52d52",
  2378 => x"5271712e",
  2379 => x"87388151",
  2380 => x"80cabd04",
  2381 => x"81135380",
  2382 => x"ca920480",
  2383 => x"517080ef",
  2384 => x"b80c0298",
  2385 => x"050d0481",
  2386 => x"0b80efb8",
  2387 => x"0c04810b",
  2388 => x"80efb80c",
  2389 => x"04810b80",
  2390 => x"efb80c04",
  2391 => x"810b80ef",
  2392 => x"b80c0402",
  2393 => x"e0050d79",
  2394 => x"7b80eef0",
  2395 => x"0887fc81",
  2396 => x"ff0680ee",
  2397 => x"f00c7184",
  2398 => x"2980eed4",
  2399 => x"05715680",
  2400 => x"eec41380",
  2401 => x"f52d8111",
  2402 => x"59575959",
  2403 => x"567480ee",
  2404 => x"c41781b7",
  2405 => x"2d7381ff",
  2406 => x"06527551",
  2407 => x"76085473",
  2408 => x"2d80efb8",
  2409 => x"085480ef",
  2410 => x"b8088025",
  2411 => x"a3387753",
  2412 => x"810b80ee",
  2413 => x"c41781b7",
  2414 => x"2d805275",
  2415 => x"51760854",
  2416 => x"732d80ef",
  2417 => x"b8085480",
  2418 => x"0b80efb8",
  2419 => x"08249738",
  2420 => x"7383fe80",
  2421 => x"0674982b",
  2422 => x"0780eef0",
  2423 => x"080780ee",
  2424 => x"f00c80cb",
  2425 => x"f00480ee",
  2426 => x"f0088807",
  2427 => x"80eef00c",
  2428 => x"80eef008",
  2429 => x"900780ee",
  2430 => x"f00c02a0",
  2431 => x"050d0402",
  2432 => x"ec050df4",
  2433 => x"90085480",
  2434 => x"eec00874",
  2435 => x"2e838038",
  2436 => x"7381a00a",
  2437 => x"06537280",
  2438 => x"2ebc3873",
  2439 => x"fc800a06",
  2440 => x"7081e6fc",
  2441 => x"0c749a2a",
  2442 => x"70810651",
  2443 => x"54557280",
  2444 => x"2e893874",
  2445 => x"810a0781",
  2446 => x"e6fc0c73",
  2447 => x"882a7080",
  2448 => x"ff065153",
  2449 => x"7280eebc",
  2450 => x"0b81b72d",
  2451 => x"80eec808",
  2452 => x"810580ee",
  2453 => x"c80c7380",
  2454 => x"d00a0653",
  2455 => x"72802ebc",
  2456 => x"3873fc80",
  2457 => x"0a067081",
  2458 => x"e7800c74",
  2459 => x"9b2a7081",
  2460 => x"06515455",
  2461 => x"72802e89",
  2462 => x"3874810a",
  2463 => x"0781e780",
  2464 => x"0c73882a",
  2465 => x"7080ff06",
  2466 => x"51537280",
  2467 => x"eebd0b81",
  2468 => x"b72d80ee",
  2469 => x"c8088105",
  2470 => x"80eec80c",
  2471 => x"73972a70",
  2472 => x"81065153",
  2473 => x"72802e8f",
  2474 => x"3880eef0",
  2475 => x"08e00670",
  2476 => x"80eef00c",
  2477 => x"f4900c73",
  2478 => x"9c2a7081",
  2479 => x"06515372",
  2480 => x"802e8d38",
  2481 => x"73962a81",
  2482 => x"06528051",
  2483 => x"80cae32d",
  2484 => x"739e2a70",
  2485 => x"81065153",
  2486 => x"72802e80",
  2487 => x"c3387388",
  2488 => x"2a80ff06",
  2489 => x"70535580",
  2490 => x"5180eecc",
  2491 => x"0853722d",
  2492 => x"80eef008",
  2493 => x"5380efb8",
  2494 => x"08802e9d",
  2495 => x"387480ee",
  2496 => x"bc0b81b7",
  2497 => x"2d800b80",
  2498 => x"eec40b81",
  2499 => x"b72d7281",
  2500 => x"0780eef0",
  2501 => x"0c80cea0",
  2502 => x"04728907",
  2503 => x"80eef00c",
  2504 => x"739d2a70",
  2505 => x"81065153",
  2506 => x"72802e8d",
  2507 => x"3873962a",
  2508 => x"81065281",
  2509 => x"5180cae3",
  2510 => x"2d738025",
  2511 => x"80c53873",
  2512 => x"882a7080",
  2513 => x"ff065153",
  2514 => x"7280eebd",
  2515 => x"0b81b72d",
  2516 => x"72528151",
  2517 => x"80eed008",
  2518 => x"53722d80",
  2519 => x"eef00853",
  2520 => x"80efb808",
  2521 => x"802e9538",
  2522 => x"800b80ee",
  2523 => x"c50b81b7",
  2524 => x"2d728207",
  2525 => x"80eef00c",
  2526 => x"80cf8304",
  2527 => x"728a0780",
  2528 => x"eef00c73",
  2529 => x"80eec00c",
  2530 => x"80eef008",
  2531 => x"f4900c02",
  2532 => x"94050d04",
  2533 => x"02c0050d",
  2534 => x"6170822b",
  2535 => x"81e6fc11",
  2536 => x"70085b5b",
  2537 => x"5c5e77ff",
  2538 => x"2e82a738",
  2539 => x"81e6f81e",
  2540 => x"80f52d57",
  2541 => x"769238ff",
  2542 => x"790c80ee",
  2543 => x"f0089807",
  2544 => x"80eef00c",
  2545 => x"80d1d204",
  2546 => x"77882a80",
  2547 => x"ff067881",
  2548 => x"ff06798f",
  2549 => x"2a7081ff",
  2550 => x"065f595b",
  2551 => x"5d778025",
  2552 => x"80f03881",
  2553 => x"e7841e80",
  2554 => x"f52d705a",
  2555 => x"5776802e",
  2556 => x"973880ee",
  2557 => x"f008fe80",
  2558 => x"0a067a98",
  2559 => x"2b079c07",
  2560 => x"80eef00c",
  2561 => x"80d1c704",
  2562 => x"f4940857",
  2563 => x"7681e788",
  2564 => x"1a81b72d",
  2565 => x"84800bf4",
  2566 => x"940c800b",
  2567 => x"f4940c81",
  2568 => x"195983ff",
  2569 => x"7925e138",
  2570 => x"81e78855",
  2571 => x"79547c53",
  2572 => x"7b527d51",
  2573 => x"80eedc1b",
  2574 => x"0857762d",
  2575 => x"80eef008",
  2576 => x"fe800a06",
  2577 => x"7a982b07",
  2578 => x"900780ee",
  2579 => x"f00c80d1",
  2580 => x"c7040280",
  2581 => x"c005f805",
  2582 => x"5681e788",
  2583 => x"5579547c",
  2584 => x"537b527d",
  2585 => x"5180eee4",
  2586 => x"1b085776",
  2587 => x"2d80efb8",
  2588 => x"08802e80",
  2589 => x"c8388059",
  2590 => x"81e78819",
  2591 => x"7080f52d",
  2592 => x"828007f4",
  2593 => x"940c7080",
  2594 => x"f52df494",
  2595 => x"0c578119",
  2596 => x"5983ff79",
  2597 => x"25e23880",
  2598 => x"eef00890",
  2599 => x"0787fc81",
  2600 => x"ff060284",
  2601 => x"05b90580",
  2602 => x"f52d7088",
  2603 => x"2b7c982b",
  2604 => x"07720780",
  2605 => x"eef00c5a",
  2606 => x"5880d1c7",
  2607 => x"0480eef0",
  2608 => x"08980780",
  2609 => x"eef00c7d",
  2610 => x"842981e6",
  2611 => x"fc0557ff",
  2612 => x"770c0280",
  2613 => x"c0050d04",
  2614 => x"02fc050d",
  2615 => x"80cbff2d",
  2616 => x"805180cf",
  2617 => x"942d8151",
  2618 => x"80cf942d",
  2619 => x"80eef008",
  2620 => x"f4900c02",
  2621 => x"84050d04",
  2622 => x"02f4050d",
  2623 => x"80eef408",
  2624 => x"8d8f2980",
  2625 => x"eef80805",
  2626 => x"70842980",
  2627 => x"fe800576",
  2628 => x"710c5153",
  2629 => x"80eef808",
  2630 => x"810580ee",
  2631 => x"f80c028c",
  2632 => x"050d0402",
  2633 => x"fc050d81",
  2634 => x"e7841351",
  2635 => x"028f0580",
  2636 => x"f52d7181",
  2637 => x"b72d0284",
  2638 => x"050d0402",
  2639 => x"f8050d73",
  2640 => x"51800b81",
  2641 => x"e6f81281",
  2642 => x"b72d80ee",
  2643 => x"f0085270",
  2644 => x"802e8d38",
  2645 => x"71ffbf06",
  2646 => x"80eef00c",
  2647 => x"80d2e704",
  2648 => x"71df0680",
  2649 => x"eef00c80",
  2650 => x"eef008f4",
  2651 => x"900c800b",
  2652 => x"80efb80c",
  2653 => x"0288050d",
  2654 => x"0402e805",
  2655 => x"0d777080",
  2656 => x"eef40c55",
  2657 => x"800b80ee",
  2658 => x"f80c7451",
  2659 => x"80d2bb2d",
  2660 => x"80d1f853",
  2661 => x"79527851",
  2662 => x"80c6db2d",
  2663 => x"80efb808",
  2664 => x"80efb808",
  2665 => x"555680ef",
  2666 => x"b808802e",
  2667 => x"81fd3880",
  2668 => x"efb80852",
  2669 => x"745180dd",
  2670 => x"ce2d80ef",
  2671 => x"b808802e",
  2672 => x"ad387482",
  2673 => x"2b80dd8a",
  2674 => x"0b80eee4",
  2675 => x"120c80dd",
  2676 => x"ac0b80ee",
  2677 => x"dc120c80",
  2678 => x"d99f0b80",
  2679 => x"eed4120c",
  2680 => x"80d6c40b",
  2681 => x"80eecc12",
  2682 => x"0c5480d4",
  2683 => x"d7047552",
  2684 => x"745180e5",
  2685 => x"812d7482",
  2686 => x"2b5480ef",
  2687 => x"b808802e",
  2688 => x"a93880e3",
  2689 => x"f80b80ee",
  2690 => x"e4150c80",
  2691 => x"e38e0b80",
  2692 => x"eedc150c",
  2693 => x"80e59e0b",
  2694 => x"80eed415",
  2695 => x"0c80e5c0",
  2696 => x"0b80eecc",
  2697 => x"150c80d4",
  2698 => x"d70480ca",
  2699 => x"c70b80ee",
  2700 => x"e4150c80",
  2701 => x"cace0b80",
  2702 => x"eedc150c",
  2703 => x"80cad50b",
  2704 => x"80eed415",
  2705 => x"0c80cadc",
  2706 => x"0b80eecc",
  2707 => x"150c80ef",
  2708 => x"b8085480",
  2709 => x"d5ab0481",
  2710 => x"0b81e6f8",
  2711 => x"1681b72d",
  2712 => x"74842980",
  2713 => x"eecc0580",
  2714 => x"eebc1680",
  2715 => x"f52d5375",
  2716 => x"52700851",
  2717 => x"54732d80",
  2718 => x"eef40880",
  2719 => x"eec40554",
  2720 => x"807481b7",
  2721 => x"2d80eef0",
  2722 => x"08547480",
  2723 => x"2e8d3873",
  2724 => x"80c00780",
  2725 => x"eef00c80",
  2726 => x"d5a20473",
  2727 => x"a00780ee",
  2728 => x"f00c80ee",
  2729 => x"f008f490",
  2730 => x"0c815473",
  2731 => x"80efb80c",
  2732 => x"0298050d",
  2733 => x"0402e405",
  2734 => x"0d807058",
  2735 => x"55800b81",
  2736 => x"e6f81681",
  2737 => x"b72d7482",
  2738 => x"2b53ff0b",
  2739 => x"81e6fc14",
  2740 => x"0c80fe80",
  2741 => x"17568d8e",
  2742 => x"54807670",
  2743 => x"8405580c",
  2744 => x"ff145473",
  2745 => x"8025f238",
  2746 => x"80cac70b",
  2747 => x"80eee414",
  2748 => x"0c80cace",
  2749 => x"0b80eedc",
  2750 => x"140c80ca",
  2751 => x"d50b80ee",
  2752 => x"d4140c80",
  2753 => x"cadc0b80",
  2754 => x"eecc140c",
  2755 => x"810b81e7",
  2756 => x"841681b7",
  2757 => x"2d8115b4",
  2758 => x"bc185855",
  2759 => x"817525ff",
  2760 => x"9c38800b",
  2761 => x"80eef80c",
  2762 => x"800b80ee",
  2763 => x"f40c800b",
  2764 => x"80eef00c",
  2765 => x"800b80ee",
  2766 => x"ec0c800b",
  2767 => x"f4900c02",
  2768 => x"9c050d04",
  2769 => x"02c0050d",
  2770 => x"61637184",
  2771 => x"2980ef84",
  2772 => x"0556415a",
  2773 => x"81557f74",
  2774 => x"082e82b8",
  2775 => x"3880d6e7",
  2776 => x"04805580",
  2777 => x"d9940480",
  2778 => x"0b80ef8c",
  2779 => x"1b80f52d",
  2780 => x"555c7b74",
  2781 => x"25829038",
  2782 => x"7b7c7b88",
  2783 => x"2980efa0",
  2784 => x"055f5f5f",
  2785 => x"81588060",
  2786 => x"75291d58",
  2787 => x"55747725",
  2788 => x"a0387982",
  2789 => x"2b1a7085",
  2790 => x"2b81eb88",
  2791 => x"05575474",
  2792 => x"167080f5",
  2793 => x"2d790581",
  2794 => x"17575954",
  2795 => x"767524ef",
  2796 => x"3881187d",
  2797 => x"0c80f098",
  2798 => x"52798d8f",
  2799 => x"2978812c",
  2800 => x"05708429",
  2801 => x"80fe8005",
  2802 => x"70085351",
  2803 => x"549d822d",
  2804 => x"80f09878",
  2805 => x"8106555b",
  2806 => x"73802e85",
  2807 => x"3882801b",
  2808 => x"5b8a5380",
  2809 => x"e9f0527a",
  2810 => x"5180ca86",
  2811 => x"2d80efb8",
  2812 => x"08feee38",
  2813 => x"79822b95",
  2814 => x"1c80f52d",
  2815 => x"7080efb0",
  2816 => x"130c80ef",
  2817 => x"b8085755",
  2818 => x"5780efb8",
  2819 => x"08742580",
  2820 => x"da38981b",
  2821 => x"58885377",
  2822 => x"52791770",
  2823 => x"852b7f84",
  2824 => x"2b057688",
  2825 => x"291181ed",
  2826 => x"c8055355",
  2827 => x"5980c7de",
  2828 => x"2d80ef98",
  2829 => x"17085675",
  2830 => x"a2387b1f",
  2831 => x"79822b05",
  2832 => x"7511832b",
  2833 => x"81edc811",
  2834 => x"51515475",
  2835 => x"861581b7",
  2836 => x"2d941b80",
  2837 => x"f52d8715",
  2838 => x"81b72d81",
  2839 => x"15881959",
  2840 => x"5580efb0",
  2841 => x"17087524",
  2842 => x"ffab3881",
  2843 => x"1c841e7f",
  2844 => x"85056189",
  2845 => x"0580ef8c",
  2846 => x"1e80f52d",
  2847 => x"5842405e",
  2848 => x"5c737c24",
  2849 => x"fdfe3879",
  2850 => x"842980ef",
  2851 => x"84056071",
  2852 => x"0c548155",
  2853 => x"7480efb8",
  2854 => x"0c0280c0",
  2855 => x"050d0402",
  2856 => x"ec050d76",
  2857 => x"787a7282",
  2858 => x"2b555654",
  2859 => x"55728025",
  2860 => x"8b3880ef",
  2861 => x"b0120851",
  2862 => x"80d9ee04",
  2863 => x"ff517280",
  2864 => x"efb01308",
  2865 => x"25a83873",
  2866 => x"88297410",
  2867 => x"05751382",
  2868 => x"2b710514",
  2869 => x"70882981",
  2870 => x"edc80581",
  2871 => x"1180f52d",
  2872 => x"821280f5",
  2873 => x"2d71882b",
  2874 => x"07525551",
  2875 => x"51517080",
  2876 => x"efb80c02",
  2877 => x"94050d04",
  2878 => x"02ffbc05",
  2879 => x"0d626468",
  2880 => x"6a6c0294",
  2881 => x"0580d705",
  2882 => x"80f52d42",
  2883 => x"425c4159",
  2884 => x"5c807887",
  2885 => x"2c7980ff",
  2886 => x"067e8429",
  2887 => x"80efb005",
  2888 => x"7008745f",
  2889 => x"5a575a58",
  2890 => x"5b7a7625",
  2891 => x"80d23876",
  2892 => x"84291770",
  2893 => x"90297da0",
  2894 => x"29057d81",
  2895 => x"80291181",
  2896 => x"edc80557",
  2897 => x"51548215",
  2898 => x"80f52d54",
  2899 => x"7c742e09",
  2900 => x"81068c38",
  2901 => x"811580f5",
  2902 => x"2d407760",
  2903 => x"2ea23887",
  2904 => x"1580f52d",
  2905 => x"861680f5",
  2906 => x"2d71882b",
  2907 => x"077c0581",
  2908 => x"1c881858",
  2909 => x"5c5c4175",
  2910 => x"7a24cb38",
  2911 => x"80dcfd04",
  2912 => x"79762581",
  2913 => x"f838807c",
  2914 => x"10187084",
  2915 => x"2980efa0",
  2916 => x"057d882a",
  2917 => x"71080573",
  2918 => x"5f5b5155",
  2919 => x"5d787d2e",
  2920 => x"80da3876",
  2921 => x"88297710",
  2922 => x"057c8429",
  2923 => x"1d567584",
  2924 => x"29057a11",
  2925 => x"832b81ed",
  2926 => x"c8117057",
  2927 => x"51515573",
  2928 => x"70810555",
  2929 => x"80f52d79",
  2930 => x"81b72d73",
  2931 => x"80f52d81",
  2932 => x"1a81b72d",
  2933 => x"821580f5",
  2934 => x"2d821a81",
  2935 => x"b72d8315",
  2936 => x"80f52d83",
  2937 => x"1a81b72d",
  2938 => x"841580f5",
  2939 => x"2d841a81",
  2940 => x"b72d8515",
  2941 => x"80f52d85",
  2942 => x"1a81b72d",
  2943 => x"7b8d8f29",
  2944 => x"78812a05",
  2945 => x"70842980",
  2946 => x"fe800570",
  2947 => x"08515154",
  2948 => x"7a742e8c",
  2949 => x"3880f098",
  2950 => x"5273519d",
  2951 => x"822d735b",
  2952 => x"80f09878",
  2953 => x"81065855",
  2954 => x"76802e85",
  2955 => x"38828015",
  2956 => x"557c1f82",
  2957 => x"801e811a",
  2958 => x"5a5a567d",
  2959 => x"802e9038",
  2960 => x"82805374",
  2961 => x"52755180",
  2962 => x"c7de2d80",
  2963 => x"dcee0482",
  2964 => x"80537552",
  2965 => x"745180c7",
  2966 => x"de2d7c82",
  2967 => x"802e8638",
  2968 => x"76802e8a",
  2969 => x"3880f098",
  2970 => x"5273519b",
  2971 => x"bf2d785d",
  2972 => x"83ff7925",
  2973 => x"ff863881",
  2974 => x"5480dcff",
  2975 => x"04805473",
  2976 => x"80efb80c",
  2977 => x"0280c405",
  2978 => x"0d0402e0",
  2979 => x"050d02b3",
  2980 => x"0580f52d",
  2981 => x"5881577e",
  2982 => x"567d5577",
  2983 => x"547b537a",
  2984 => x"52795180",
  2985 => x"d9f82d02",
  2986 => x"a0050d04",
  2987 => x"02e0050d",
  2988 => x"02b30580",
  2989 => x"f52d5880",
  2990 => x"5780567d",
  2991 => x"5577547b",
  2992 => x"537a5279",
  2993 => x"5180d9f8",
  2994 => x"2d02a005",
  2995 => x"0d0402d8",
  2996 => x"050d7b80",
  2997 => x"f0985370",
  2998 => x"b4bc2980",
  2999 => x"fe800570",
  3000 => x"08535559",
  3001 => x"9d822d88",
  3002 => x"5380f098",
  3003 => x"5280eacc",
  3004 => x"5180ca86",
  3005 => x"2d80efb8",
  3006 => x"0880fa38",
  3007 => x"78822b56",
  3008 => x"810b80ef",
  3009 => x"98170c80",
  3010 => x"f0c80b80",
  3011 => x"f52d7080",
  3012 => x"ef90180c",
  3013 => x"5580f0c9",
  3014 => x"0b80f52d",
  3015 => x"80ef8c1a",
  3016 => x"81b72d80",
  3017 => x"efb80854",
  3018 => x"7480d024",
  3019 => x"81e33880",
  3020 => x"efb80880",
  3021 => x"ef8c1a80",
  3022 => x"f52d7671",
  3023 => x"29565957",
  3024 => x"80efb808",
  3025 => x"742581bc",
  3026 => x"38781685",
  3027 => x"2b81eb88",
  3028 => x"05757929",
  3029 => x"80f0cc5a",
  3030 => x"56567616",
  3031 => x"54777081",
  3032 => x"055980f5",
  3033 => x"2d7481b7",
  3034 => x"2d811757",
  3035 => x"747724ea",
  3036 => x"3880e084",
  3037 => x"04885380",
  3038 => x"f0985280",
  3039 => x"eac05180",
  3040 => x"ca862d80",
  3041 => x"5480efb8",
  3042 => x"08742e09",
  3043 => x"81068181",
  3044 => x"3878822b",
  3045 => x"80f0c80b",
  3046 => x"80f52d70",
  3047 => x"80ef9013",
  3048 => x"0c565680",
  3049 => x"f0c90b80",
  3050 => x"f52d80ef",
  3051 => x"8c1a81b7",
  3052 => x"2d80efb8",
  3053 => x"0880ef98",
  3054 => x"170c80ef",
  3055 => x"b8085474",
  3056 => x"80d02480",
  3057 => x"cc3880ef",
  3058 => x"b80880ef",
  3059 => x"8c1a80f5",
  3060 => x"2d767129",
  3061 => x"56595780",
  3062 => x"efb80874",
  3063 => x"25a63878",
  3064 => x"16852b81",
  3065 => x"eb880575",
  3066 => x"792980f0",
  3067 => x"cb0b80f5",
  3068 => x"2d57575a",
  3069 => x"761a5474",
  3070 => x"7481b72d",
  3071 => x"81175775",
  3072 => x"7724f138",
  3073 => x"78842980",
  3074 => x"ef840554",
  3075 => x"ff740c81",
  3076 => x"547380ef",
  3077 => x"b80c02a8",
  3078 => x"050d0402",
  3079 => x"e8050d77",
  3080 => x"7957548c",
  3081 => x"5380eab0",
  3082 => x"52735180",
  3083 => x"c7de2d75",
  3084 => x"901581b7",
  3085 => x"2d800b91",
  3086 => x"1581b72d",
  3087 => x"820b9415",
  3088 => x"81b72d89",
  3089 => x"0b951581",
  3090 => x"b72d80d2",
  3091 => x"0b961581",
  3092 => x"b72de50b",
  3093 => x"971581b7",
  3094 => x"2d805575",
  3095 => x"981581b7",
  3096 => x"2d800b99",
  3097 => x"1581b72d",
  3098 => x"80eaa415",
  3099 => x"80f52d9a",
  3100 => x"1581b72d",
  3101 => x"820b9b15",
  3102 => x"81b72d82",
  3103 => x"0b9f1581",
  3104 => x"b72d8115",
  3105 => x"88155555",
  3106 => x"887525cf",
  3107 => x"38029805",
  3108 => x"0d0402e8",
  3109 => x"050d7780",
  3110 => x"eefc0856",
  3111 => x"54815674",
  3112 => x"80cd3884",
  3113 => x"80537452",
  3114 => x"735180c8",
  3115 => x"892da553",
  3116 => x"80e9fc52",
  3117 => x"735180c7",
  3118 => x"de2da80b",
  3119 => x"b01581b7",
  3120 => x"2d810bb1",
  3121 => x"1581b72d",
  3122 => x"a8539352",
  3123 => x"b4145180",
  3124 => x"c8892d74",
  3125 => x"52828014",
  3126 => x"5180e09b",
  3127 => x"2d80eefc",
  3128 => x"081680ee",
  3129 => x"fc0c7480",
  3130 => x"ef800c80",
  3131 => x"e2c70480",
  3132 => x"ef800881",
  3133 => x"0580ef80",
  3134 => x"0c80ef80",
  3135 => x"08932e09",
  3136 => x"8106ab38",
  3137 => x"82805380",
  3138 => x"52735180",
  3139 => x"c8892d80",
  3140 => x"eefc0852",
  3141 => x"80eefc08",
  3142 => x"810580ee",
  3143 => x"fc0c7351",
  3144 => x"80e09b2d",
  3145 => x"800b80ef",
  3146 => x"800c80e2",
  3147 => x"ba048280",
  3148 => x"5381e552",
  3149 => x"735180c8",
  3150 => x"892d8280",
  3151 => x"14ff1757",
  3152 => x"54758025",
  3153 => x"ffa93881",
  3154 => x"0b80efb8",
  3155 => x"0c029805",
  3156 => x"0d0402f4",
  3157 => x"050d800b",
  3158 => x"80eefc0c",
  3159 => x"8bf28053",
  3160 => x"80e19252",
  3161 => x"745180c5",
  3162 => x"a92d028c",
  3163 => x"050d0402",
  3164 => x"f8050d74",
  3165 => x"84291576",
  3166 => x"88291771",
  3167 => x"88290578",
  3168 => x"05febf05",
  3169 => x"80efb80c",
  3170 => x"51028805",
  3171 => x"0d0402e4",
  3172 => x"050d7802",
  3173 => x"8405af05",
  3174 => x"80f52d55",
  3175 => x"7b547a53",
  3176 => x"70525780",
  3177 => x"e2ef2d80",
  3178 => x"5680efb8",
  3179 => x"088d8e26",
  3180 => x"bd38768d",
  3181 => x"8f2980ef",
  3182 => x"b8080570",
  3183 => x"842980fe",
  3184 => x"80057008",
  3185 => x"515155bd",
  3186 => x"b12d7480",
  3187 => x"efb80827",
  3188 => x"9d38bdb1",
  3189 => x"2d7480ef",
  3190 => x"b8082792",
  3191 => x"387c5274",
  3192 => x"519bbf2d",
  3193 => x"80efb808",
  3194 => x"762e8338",
  3195 => x"81567580",
  3196 => x"efb80c02",
  3197 => x"9c050d04",
  3198 => x"02d4050d",
  3199 => x"7c7e6064",
  3200 => x"029005bf",
  3201 => x"0580f52d",
  3202 => x"70597258",
  3203 => x"73577456",
  3204 => x"5c5a5c5c",
  3205 => x"5980e2ef",
  3206 => x"2d805680",
  3207 => x"efb8088d",
  3208 => x"8e2680d3",
  3209 => x"38788d8f",
  3210 => x"2980efb8",
  3211 => x"08057084",
  3212 => x"2980fe80",
  3213 => x"05700851",
  3214 => x"5155bdb1",
  3215 => x"2d7480ef",
  3216 => x"b80827b3",
  3217 => x"38797781",
  3218 => x"b72d7a81",
  3219 => x"1881b72d",
  3220 => x"77821881",
  3221 => x"b72d820b",
  3222 => x"831881b7",
  3223 => x"2d800b84",
  3224 => x"1881b72d",
  3225 => x"800b8518",
  3226 => x"81b72d60",
  3227 => x"5274519d",
  3228 => x"822d80ef",
  3229 => x"b8085675",
  3230 => x"80efb80c",
  3231 => x"02ac050d",
  3232 => x"0402f805",
  3233 => x"0d748ba0",
  3234 => x"80327009",
  3235 => x"81057072",
  3236 => x"07802580",
  3237 => x"efb80c52",
  3238 => x"52028805",
  3239 => x"0d0402f8",
  3240 => x"050d7451",
  3241 => x"89528071",
  3242 => x"248c3881",
  3243 => x"c1115288",
  3244 => x"71258338",
  3245 => x"ff527180",
  3246 => x"efb80c02",
  3247 => x"88050d04",
  3248 => x"810b80ef",
  3249 => x"b80c0400",
  3250 => x"00ffffff",
  3251 => x"ff00ffff",
  3252 => x"ffff00ff",
  3253 => x"ffffff00",
  3254 => x"000055aa",
  3255 => x"00000000",
  3256 => x"496e7365",
  3257 => x"72742064",
  3258 => x"69736b20",
  3259 => x"30000000",
  3260 => x"57726974",
  3261 => x"65207072",
  3262 => x"6f746563",
  3263 => x"74206469",
  3264 => x"736b2030",
  3265 => x"00000000",
  3266 => x"496e7365",
  3267 => x"72742064",
  3268 => x"69736b20",
  3269 => x"31000000",
  3270 => x"57726974",
  3271 => x"65207072",
  3272 => x"6f746563",
  3273 => x"74206469",
  3274 => x"736b2031",
  3275 => x"00000000",
  3276 => x"43726561",
  3277 => x"74652062",
  3278 => x"6c616e6b",
  3279 => x"20646973",
  3280 => x"6b000000",
  3281 => x"4261636b",
  3282 => x"00000000",
  3283 => x"4469736b",
  3284 => x"206d656e",
  3285 => x"75202020",
  3286 => x"20202020",
  3287 => x"20202020",
  3288 => x"20100000",
  3289 => x"45786974",
  3290 => x"00000000",
  3291 => x"4469736b",
  3292 => x"206d656e",
  3293 => x"752e0000",
  3294 => x"4c6f6164",
  3295 => x"696e6720",
  3296 => x"6661696c",
  3297 => x"65640000",
  3298 => x"4f4b0000",
  3299 => x"4c6f6164",
  3300 => x"696e6720",
  3301 => x"524f4d73",
  3302 => x"2e2e2e0a",
  3303 => x"2e2e2e66",
  3304 => x"726f6d20",
  3305 => x"2f414d53",
  3306 => x"54524144",
  3307 => x"2f414d53",
  3308 => x"444f532e",
  3309 => x"524f4d2e",
  3310 => x"2e2e0000",
  3311 => x"414d5354",
  3312 => x"52414400",
  3313 => x"414d5344",
  3314 => x"4f532e52",
  3315 => x"4f4d0000",
  3316 => x"42415349",
  3317 => x"43312d31",
  3318 => x"2e524f4d",
  3319 => x"00000000",
  3320 => x"4661696c",
  3321 => x"65642074",
  3322 => x"6f206368",
  3323 => x"616e6765",
  3324 => x"20646972",
  3325 => x"6563746f",
  3326 => x"72790000",
  3327 => x"4449534b",
  3328 => x"00000000",
  3329 => x"2e494d47",
  3330 => x"00000000",
  3331 => x"43726561",
  3332 => x"74696e67",
  3333 => x"2066696c",
  3334 => x"653a2000",
  3335 => x"496e6974",
  3336 => x"69616c69",
  3337 => x"7a696e67",
  3338 => x"20534420",
  3339 => x"63617264",
  3340 => x"0a000000",
  3341 => x"14200000",
  3342 => x"15200000",
  3343 => x"53442069",
  3344 => x"6e69742e",
  3345 => x"2e2e0a00",
  3346 => x"53442063",
  3347 => x"61726420",
  3348 => x"72657365",
  3349 => x"74206661",
  3350 => x"696c6564",
  3351 => x"210a0000",
  3352 => x"53444843",
  3353 => x"20657272",
  3354 => x"6f72210a",
  3355 => x"00000000",
  3356 => x"57726974",
  3357 => x"65206661",
  3358 => x"696c6564",
  3359 => x"0a000000",
  3360 => x"52656164",
  3361 => x"20666169",
  3362 => x"6c65640a",
  3363 => x"00000000",
  3364 => x"43617264",
  3365 => x"20696e69",
  3366 => x"74206661",
  3367 => x"696c6564",
  3368 => x"0a000000",
  3369 => x"46415431",
  3370 => x"36202020",
  3371 => x"00000000",
  3372 => x"46415433",
  3373 => x"32202020",
  3374 => x"00000000",
  3375 => x"4e6f2070",
  3376 => x"61727469",
  3377 => x"74696f6e",
  3378 => x"20736967",
  3379 => x"0a000000",
  3380 => x"42616420",
  3381 => x"70617274",
  3382 => x"0a000000",
  3383 => x"30313233",
  3384 => x"34353637",
  3385 => x"38396162",
  3386 => x"63646566",
  3387 => x"00000000",
  3388 => x"54726163",
  3389 => x"6b2d496e",
  3390 => x"666f0000",
  3391 => x"45585445",
  3392 => x"4e444544",
  3393 => x"20446973",
  3394 => x"6b2d4669",
  3395 => x"6c650d0a",
  3396 => x"43504345",
  3397 => x"43203230",
  3398 => x"32323034",
  3399 => x"31320d0a",
  3400 => x"1a000000",
  3401 => x"c1c6c2c7",
  3402 => x"c3c8c4c9",
  3403 => x"c5000000",
  3404 => x"54726163",
  3405 => x"6b2d496e",
  3406 => x"666f0d0a",
  3407 => x"00000000",
  3408 => x"4d56202d",
  3409 => x"20435043",
  3410 => x"00000000",
  3411 => x"45585445",
  3412 => x"4e444544",
  3413 => x"00000000",
  3414 => x"00000002",
  3415 => x"00000004",
  3416 => x"0000334c",
  3417 => x"00003580",
  3418 => x"00000002",
  3419 => x"00003364",
  3420 => x"000007c1",
  3421 => x"00000000",
  3422 => x"00000000",
  3423 => x"00000000",
  3424 => x"00000004",
  3425 => x"0000336c",
  3426 => x"00003580",
  3427 => x"00000004",
  3428 => x"0000346c",
  3429 => x"00003580",
  3430 => x"00000002",
  3431 => x"000032e0",
  3432 => x"000003b2",
  3433 => x"00000001",
  3434 => x"000032f0",
  3435 => x"00000006",
  3436 => x"00000002",
  3437 => x"00003308",
  3438 => x"000003d1",
  3439 => x"00000001",
  3440 => x"00003318",
  3441 => x"00000007",
  3442 => x"00000002",
  3443 => x"00003330",
  3444 => x"000003f0",
  3445 => x"00000004",
  3446 => x"0000346c",
  3447 => x"00003580",
  3448 => x"00000004",
  3449 => x"00003344",
  3450 => x"0000355c",
  3451 => x"00000000",
  3452 => x"00000000",
  3453 => x"00000000",
  3454 => x"00000004",
  3455 => x"00003378",
  3456 => x"000035f8",
  3457 => x"00000004",
  3458 => x"00003388",
  3459 => x"0000355c",
  3460 => x"00000000",
  3461 => x"00000000",
  3462 => x"00000000",
  3463 => x"00000000",
  3464 => x"00000000",
  3465 => x"00000000",
  3466 => x"00000000",
  3467 => x"00000000",
  3468 => x"00000000",
  3469 => x"00000000",
  3470 => x"00000000",
  3471 => x"00000000",
  3472 => x"00000000",
  3473 => x"00000000",
  3474 => x"00000000",
  3475 => x"00000000",
  3476 => x"00000000",
  3477 => x"00000000",
  3478 => x"00000000",
  3479 => x"00000000",
  3480 => x"00000000",
  3481 => x"00000000",
  3482 => x"00000000",
  3483 => x"00000000",
  3484 => x"000000c6",
  3485 => x"00000000",
  3486 => x"00000000",
  3487 => x"7fffffff",
  3488 => x"00000002",
  3489 => x"00000002",
  3490 => x"00003d6c",
  3491 => x"0000205d",
  3492 => x"00000002",
  3493 => x"00003d8a",
  3494 => x"0000205d",
  3495 => x"00000002",
  3496 => x"00003da8",
  3497 => x"0000205d",
  3498 => x"00000002",
  3499 => x"00003dc6",
  3500 => x"0000205d",
  3501 => x"00000002",
  3502 => x"00003de4",
  3503 => x"0000205d",
  3504 => x"00000002",
  3505 => x"00003e02",
  3506 => x"0000205d",
  3507 => x"00000002",
  3508 => x"00003e20",
  3509 => x"0000205d",
  3510 => x"00000002",
  3511 => x"00003e3e",
  3512 => x"0000205d",
  3513 => x"00000002",
  3514 => x"00003e5c",
  3515 => x"0000205d",
  3516 => x"00000002",
  3517 => x"00003e7a",
  3518 => x"0000205d",
  3519 => x"00000002",
  3520 => x"00003e98",
  3521 => x"0000205d",
  3522 => x"00000002",
  3523 => x"00003eb6",
  3524 => x"0000205d",
  3525 => x"00000002",
  3526 => x"00003ed4",
  3527 => x"0000205d",
  3528 => x"00000004",
  3529 => x"00003344",
  3530 => x"00000000",
  3531 => x"00000000",
  3532 => x"00000000",
  3533 => x"000020e3",
  3534 => x"00000000",
  3535 => x"00000000",
  3536 => x"00000000",
  3537 => x"00000000",
  3538 => x"00000000",
  3539 => x"00000000",
  3540 => x"00000000",
  3541 => x"00000000",
  3542 => x"00000000",
  3543 => x"00000000",
  3544 => x"00000000",
  3545 => x"00000000",
  3546 => x"00000000",
  3547 => x"00000000",
  3548 => x"00000000",
  3549 => x"00000000",
  3550 => x"00000000",
  3551 => x"00000000",
  3552 => x"00000000",
  3553 => x"ffffffff",
  3554 => x"00000000",
  3555 => x"00000000",
  3556 => x"00000000",
  3557 => x"00000000",
  3558 => x"00000000",
  3559 => x"00000000",
  3560 => x"00000000",
  3561 => x"00000000",
  3562 => x"00000000",
  3563 => x"00000000",
  3564 => x"00000000",
  3565 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

